# 
# LEF OUT 
# User Name : bcruik2 
# Date : Sat Mar 21 12:22:37 2020
# 
VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MANUFACTURINGGRID 0.001 ;

LAYER NWELL
  TYPE MASTERSLICE ;
END NWELL

LAYER DNW
  TYPE MASTERSLICE ;
END DNW

LAYER DIFF
  TYPE MASTERSLICE ;
END DIFF

LAYER PIMP
  TYPE MASTERSLICE ;
END PIMP

LAYER NIMP
  TYPE MASTERSLICE ;
END NIMP

LAYER DIFF_18
  TYPE MASTERSLICE ;
END DIFF_18

LAYER PAD
  TYPE MASTERSLICE ;
END PAD

LAYER ESD_25
  TYPE MASTERSLICE ;
END ESD_25

LAYER SBLK
  TYPE MASTERSLICE ;
END SBLK

LAYER HVTIMP
  TYPE MASTERSLICE ;
END HVTIMP

LAYER LVTIMP
  TYPE MASTERSLICE ;
END LVTIMP

LAYER M1PIN
  TYPE MASTERSLICE ;
END M1PIN

LAYER M2PIN
  TYPE MASTERSLICE ;
END M2PIN

LAYER M3PIN
  TYPE MASTERSLICE ;
END M3PIN

LAYER M4PIN
  TYPE MASTERSLICE ;
END M4PIN

LAYER M5PIN
  TYPE MASTERSLICE ;
END M5PIN

LAYER M6PIN
  TYPE MASTERSLICE ;
END M6PIN

LAYER M7PIN
  TYPE MASTERSLICE ;
END M7PIN

LAYER M8PIN
  TYPE MASTERSLICE ;
END M8PIN

LAYER M9PIN
  TYPE MASTERSLICE ;
END M9PIN

LAYER MRDL9PIN
  TYPE MASTERSLICE ;
END MRDL9PIN

LAYER HOTNWL
  TYPE MASTERSLICE ;
END HOTNWL

LAYER DIOD
  TYPE MASTERSLICE ;
END DIOD

LAYER BJTDMY
  TYPE MASTERSLICE ;
END BJTDMY

LAYER RNW
  TYPE MASTERSLICE ;
END RNW

LAYER RMARK
  TYPE MASTERSLICE ;
END RMARK

LAYER prBoundary
  TYPE MASTERSLICE ;
END prBoundary

LAYER LOGO
  TYPE MASTERSLICE ;
END LOGO

LAYER IP
  TYPE MASTERSLICE ;
END IP

LAYER RM1
  TYPE MASTERSLICE ;
END RM1

LAYER RM2
  TYPE MASTERSLICE ;
END RM2

LAYER RM3
  TYPE MASTERSLICE ;
END RM3

LAYER RM4
  TYPE MASTERSLICE ;
END RM4

LAYER RM5
  TYPE MASTERSLICE ;
END RM5

LAYER RM6
  TYPE MASTERSLICE ;
END RM6

LAYER RM7
  TYPE MASTERSLICE ;
END RM7

LAYER RM8
  TYPE MASTERSLICE ;
END RM8

LAYER RM9
  TYPE MASTERSLICE ;
END RM9

LAYER DM1EXCL
  TYPE MASTERSLICE ;
END DM1EXCL

LAYER DM2EXCL
  TYPE MASTERSLICE ;
END DM2EXCL

LAYER DM3EXCL
  TYPE MASTERSLICE ;
END DM3EXCL

LAYER DM4EXCL
  TYPE MASTERSLICE ;
END DM4EXCL

LAYER DM5EXCL
  TYPE MASTERSLICE ;
END DM5EXCL

LAYER DM6EXCL
  TYPE MASTERSLICE ;
END DM6EXCL

LAYER DM7EXCL
  TYPE MASTERSLICE ;
END DM7EXCL

LAYER DM8EXCL
  TYPE MASTERSLICE ;
END DM8EXCL

LAYER DM9EXCL
  TYPE MASTERSLICE ;
END DM9EXCL

LAYER DIFF_25
  TYPE MASTERSLICE ;
END DIFF_25

LAYER DIFF_FM
  TYPE MASTERSLICE ;
END DIFF_FM

LAYER PO_FM
  TYPE MASTERSLICE ;
END PO_FM

LAYER PO
  TYPE MASTERSLICE ;
END PO

LAYER CO
  TYPE CUT ;
  SPACING 0.05 ;
END CO

LAYER M1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.152 ;
  WIDTH 0.05 ;
  AREA 0.01 ;
  MAXWIDTH 5 ;
  MINWIDTH 0.05 ;
  SPACING 0.05 ;
  MINENCLOSEDAREA 0.2 ;
  CAPMULTIPLIER 1 ;
  PROTRUSIONWIDTH 0.06 LENGTH 0.1 WIDTH 0.15 ;
  PROTRUSIONWIDTH 0.07 LENGTH 0.17 WIDTH 0.3 ;
  PROTRUSIONWIDTH 0.15 LENGTH 0.7 WIDTH 1.5 ;
  MINIMUMDENSITY 10 ;
  MAXIMUMDENSITY 85 ;
  DENSITYCHECKWINDOW 75 75 ;
  DENSITYCHECKSTEP 37.5 ;
  MINIMUMDENSITY 1 ;
  MAXIMUMDENSITY 60 ;
  DENSITYCHECKWINDOW 100 100 ;
  DENSITYCHECKSTEP 50 ;
END M1

LAYER VIA1
  TYPE CUT ;
  SPACING 0.07 ;
END VIA1

LAYER M2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.152 ;
  WIDTH 0.056 ;
  AREA 0.016 ;
  MAXWIDTH 5 ;
  MINWIDTH 0.056 ;
  SPACING 0.056 ;
  MINENCLOSEDAREA 0.2 ;
  CAPMULTIPLIER 1 ;
  PROTRUSIONWIDTH 0.06 LENGTH 0.1 WIDTH 0.15 ;
  PROTRUSIONWIDTH 0.07 LENGTH 0.15 WIDTH 0.3 ;
  PROTRUSIONWIDTH 0.15 LENGTH 0.7 WIDTH 1.5 ;
  PROTRUSIONWIDTH 0.3 LENGTH 1.5 WIDTH 3 ;
  MINIMUMDENSITY 15 ;
  MAXIMUMDENSITY 100 ;
  DENSITYCHECKWINDOW 50 50 ;
  DENSITYCHECKSTEP 25 ;
  MINIMUMDENSITY 1 ;
  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 100 100 ;
  DENSITYCHECKSTEP 50 ;
END M2

LAYER VIA2
  TYPE CUT ;
  SPACING 0.07 ;
END VIA2

LAYER M3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.304 ;
  WIDTH 0.056 ;
  AREA 0.016 ;
  MAXWIDTH 5 ;
  MINWIDTH 0.056 ;
  SPACING 0.056 ;
  MINENCLOSEDAREA 0.2 ;
  CAPMULTIPLIER 1 ;
  PROTRUSIONWIDTH 0.06 LENGTH 0.1 WIDTH 0.15 ;
  PROTRUSIONWIDTH 0.07 LENGTH 0.15 WIDTH 0.3 ;
  PROTRUSIONWIDTH 0.15 LENGTH 0.7 WIDTH 1.5 ;
  PROTRUSIONWIDTH 0.3 LENGTH 1.5 WIDTH 3 ;
  MINIMUMDENSITY 15 ;
  MAXIMUMDENSITY 100 ;
  DENSITYCHECKWINDOW 50 50 ;
  DENSITYCHECKSTEP 25 ;
  MINIMUMDENSITY 1 ;
  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 100 100 ;
  DENSITYCHECKSTEP 50 ;
END M3

LAYER VIA3
  TYPE CUT ;
  SPACING 0.07 ;
END VIA3

LAYER M4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.304 ;
  WIDTH 0.056 ;
  AREA 0.016 ;
  MAXWIDTH 5 ;
  MINWIDTH 0.056 ;
  SPACING 0.056 ;
  MINENCLOSEDAREA 0.2 ;
  CAPMULTIPLIER 1 ;
  PROTRUSIONWIDTH 0.06 LENGTH 0.1 WIDTH 0.15 ;
  PROTRUSIONWIDTH 0.07 LENGTH 0.15 WIDTH 0.3 ;
  PROTRUSIONWIDTH 0.15 LENGTH 0.7 WIDTH 1.5 ;
  PROTRUSIONWIDTH 0.3 LENGTH 1.5 WIDTH 3 ;
  MINIMUMDENSITY 15 ;
  MAXIMUMDENSITY 100 ;
  DENSITYCHECKWINDOW 50 50 ;
  DENSITYCHECKSTEP 25 ;
  MINIMUMDENSITY 1 ;
  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 100 100 ;
  DENSITYCHECKSTEP 50 ;
END M4

LAYER VIA4
  TYPE CUT ;
  SPACING 0.07 ;
END VIA4

LAYER M5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.608 ;
  WIDTH 0.056 ;
  AREA 0.016 ;
  MAXWIDTH 5 ;
  MINWIDTH 0.056 ;
  SPACING 0.056 ;
  MINENCLOSEDAREA 0.2 ;
  CAPMULTIPLIER 1 ;
  PROTRUSIONWIDTH 0.06 LENGTH 0.1 WIDTH 0.15 ;
  PROTRUSIONWIDTH 0.07 LENGTH 0.15 WIDTH 0.3 ;
  PROTRUSIONWIDTH 0.15 LENGTH 0.7 WIDTH 1.5 ;
  PROTRUSIONWIDTH 0.3 LENGTH 1.5 WIDTH 3 ;
  MINIMUMDENSITY 15 ;
  MAXIMUMDENSITY 100 ;
  DENSITYCHECKWINDOW 50 50 ;
  DENSITYCHECKSTEP 25 ;
  MINIMUMDENSITY 1 ;
  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 100 100 ;
  DENSITYCHECKSTEP 50 ;
END M5

LAYER VIA5
  TYPE CUT ;
  SPACING 0.07 ;
END VIA5

LAYER M6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.608 ;
  WIDTH 0.056 ;
  AREA 0.016 ;
  MAXWIDTH 5 ;
  MINWIDTH 0.056 ;
  SPACING 0.056 ;
  MINENCLOSEDAREA 0.2 ;
  CAPMULTIPLIER 1 ;
  PROTRUSIONWIDTH 0.06 LENGTH 0.1 WIDTH 0.15 ;
  PROTRUSIONWIDTH 0.07 LENGTH 0.15 WIDTH 0.3 ;
  PROTRUSIONWIDTH 0.15 LENGTH 0.7 WIDTH 1.5 ;
  PROTRUSIONWIDTH 0.3 LENGTH 1.5 WIDTH 3 ;
  MINIMUMDENSITY 15 ;
  MAXIMUMDENSITY 100 ;
  DENSITYCHECKWINDOW 50 50 ;
  DENSITYCHECKSTEP 25 ;
  MINIMUMDENSITY 1 ;
  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 100 100 ;
  DENSITYCHECKSTEP 50 ;
END M6

LAYER VIA6
  TYPE CUT ;
  SPACING 0.07 ;
END VIA6

LAYER M7
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 1.216 ;
  WIDTH 0.056 ;
  AREA 0.016 ;
  MAXWIDTH 5 ;
  MINWIDTH 0.056 ;
  SPACING 0.056 ;
  MINENCLOSEDAREA 0.2 ;
  CAPMULTIPLIER 1 ;
  PROTRUSIONWIDTH 0.06 LENGTH 0.1 WIDTH 0.15 ;
  PROTRUSIONWIDTH 0.07 LENGTH 0.15 WIDTH 0.3 ;
  PROTRUSIONWIDTH 0.15 LENGTH 0.7 WIDTH 1.5 ;
  PROTRUSIONWIDTH 0.3 LENGTH 1.5 WIDTH 3 ;
  MINIMUMDENSITY 15 ;
  MAXIMUMDENSITY 100 ;
  DENSITYCHECKWINDOW 50 50 ;
  DENSITYCHECKSTEP 25 ;
  MINIMUMDENSITY 1 ;
  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 100 100 ;
  DENSITYCHECKSTEP 50 ;
END M7

LAYER VIA7
  TYPE CUT ;
  SPACING 0.07 ;
END VIA7

LAYER M8
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 1.216 ;
  WIDTH 0.056 ;
  AREA 0.016 ;
  MAXWIDTH 5 ;
  MINWIDTH 0.056 ;
  SPACING 0.056 ;
  MINENCLOSEDAREA 0.2 ;
  CAPMULTIPLIER 1 ;
  PROTRUSIONWIDTH 0.06 LENGTH 0.1 WIDTH 0.15 ;
  PROTRUSIONWIDTH 0.07 LENGTH 0.15 WIDTH 0.3 ;
  PROTRUSIONWIDTH 0.15 LENGTH 0.7 WIDTH 1.5 ;
  PROTRUSIONWIDTH 0.3 LENGTH 1.5 WIDTH 3 ;
  MINIMUMDENSITY 15 ;
  MAXIMUMDENSITY 100 ;
  DENSITYCHECKWINDOW 50 50 ;
  DENSITYCHECKSTEP 25 ;
  MINIMUMDENSITY 1 ;
  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 100 100 ;
  DENSITYCHECKSTEP 50 ;
END M8

LAYER VIA8
  TYPE CUT ;
  SPACING 0.12 ;
END VIA8

LAYER M9
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 2.432 ;
  WIDTH 0.16 ;
  AREA 0.055 ;
  MAXWIDTH 10 ;
  MINWIDTH 0.16 ;
  SPACING 0.056 ;
  MINENCLOSEDAREA 0.2 ;
  CAPMULTIPLIER 1 ;
  MINIMUMDENSITY 15 ;
  MAXIMUMDENSITY 100 ;
  DENSITYCHECKWINDOW 50 50 ;
  DENSITYCHECKSTEP 25 ;
  MINIMUMDENSITY 1 ;
  MAXIMUMDENSITY 60 ;
  DENSITYCHECKWINDOW 100 100 ;
  DENSITYCHECKSTEP 50 ;
END M9

LAYER VIARDL
  TYPE CUT ;
  SPACING 2 ;
END VIARDL

LAYER MRDL
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 4.864 ;
  WIDTH 2 ;
  AREA 4 ;
  SPACING 2 ;
  MAXWIDTH 30 ;
  MINWIDTH 2 ;
  MINENCLOSEDAREA 0.2 ;
  CAPMULTIPLIER 1 ;
END MRDL

LAYER OverlapCheck
  TYPE OVERLAP ;
END OverlapCheck

VIA VIA12SQ_C
  DEFAULT 
  RESISTANCE 1.6 ;
  LAYER M1 ;
    RECT -0.0550 -0.0300 0.0550 0.0300 ;
  LAYER VIA1 ;
    RECT -0.0250 -0.0250 0.0250 0.0250 ;
  LAYER M2 ;
    RECT -0.0300 -0.0550 0.0300 0.0550 ;
END VIA12SQ_C

VIA VIA12BAR_C
  RESISTANCE 1.6 ;
  LAYER M1 ;
    RECT -0.0550 -0.0550 0.0550 0.0550 ;
  LAYER VIA1 ;
    RECT -0.0250 -0.0500 0.0250 0.0500 ;
  LAYER M2 ;
    RECT -0.0300 -0.0800 0.0300 0.0800 ;
END VIA12BAR_C

VIA VIA12LG_C
  RESISTANCE 1.6 ;
  LAYER M1 ;
    RECT -0.0800 -0.0550 0.0800 0.0550 ;
  LAYER VIA1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0800 -0.0550 0.0800 0.0550 ;
END VIA12LG_C

VIA VIA12SQ
  RESISTANCE 1.6 ;
  LAYER M1 ;
    RECT -0.0550 -0.0300 0.0550 0.0300 ;
  LAYER VIA1 ;
    RECT -0.0250 -0.0250 0.0250 0.0250 ;
  LAYER M2 ;
    RECT -0.0550 -0.0300 0.0550 0.0300 ;
END VIA12SQ

VIA VIA12BAR
  RESISTANCE 1.6 ;
  LAYER M1 ;
    RECT -0.0550 -0.0550 0.0550 0.0550 ;
  LAYER VIA1 ;
    RECT -0.0250 -0.0500 0.0250 0.0500 ;
  LAYER M2 ;
    RECT -0.0550 -0.0550 0.0550 0.0550 ;
END VIA12BAR

VIA VIA12LG
  RESISTANCE 1.6 ;
  LAYER M1 ;
    RECT -0.0800 -0.0550 0.0800 0.0550 ;
  LAYER VIA1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M2 ;
    RECT -0.0800 -0.0550 0.0800 0.0550 ;
END VIA12LG

VIA VIA23SQ_C
  DEFAULT 
  RESISTANCE 1.6 ;
  LAYER M2 ;
    RECT -0.0550 -0.0300 0.0550 0.0300 ;
  LAYER VIA2 ;
    RECT -0.0250 -0.0250 0.0250 0.0250 ;
  LAYER M3 ;
    RECT -0.0300 -0.0550 0.0300 0.0550 ;
END VIA23SQ_C

VIA VIA23BAR_C
  RESISTANCE 1.6 ;
  LAYER M2 ;
    RECT -0.0550 -0.0550 0.0550 0.0550 ;
  LAYER VIA2 ;
    RECT -0.0250 -0.0500 0.0250 0.0500 ;
  LAYER M3 ;
    RECT -0.0300 -0.0800 0.0300 0.0800 ;
END VIA23BAR_C

VIA VIA23LG_C
  RESISTANCE 1.6 ;
  LAYER M2 ;
    RECT -0.0800 -0.0550 0.0800 0.0550 ;
  LAYER VIA2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0800 -0.0550 0.0800 0.0550 ;
END VIA23LG_C

VIA VIA23SQ
  RESISTANCE 1.6 ;
  LAYER M2 ;
    RECT -0.0550 -0.0300 0.0550 0.0300 ;
  LAYER VIA2 ;
    RECT -0.0250 -0.0250 0.0250 0.0250 ;
  LAYER M3 ;
    RECT -0.0550 -0.0300 0.0550 0.0300 ;
END VIA23SQ

VIA VIA23BAR
  RESISTANCE 1.6 ;
  LAYER M2 ;
    RECT -0.0550 -0.0550 0.0550 0.0550 ;
  LAYER VIA2 ;
    RECT -0.0250 -0.0500 0.0250 0.0500 ;
  LAYER M3 ;
    RECT -0.0550 -0.0550 0.0550 0.0550 ;
END VIA23BAR

VIA VIA23LG
  RESISTANCE 1.6 ;
  LAYER M2 ;
    RECT -0.0800 -0.0550 0.0800 0.0550 ;
  LAYER VIA2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M3 ;
    RECT -0.0800 -0.0550 0.0800 0.0550 ;
END VIA23LG

VIA VIA34SQ_C
  DEFAULT 
  RESISTANCE 1.6 ;
  LAYER M3 ;
    RECT -0.0550 -0.0300 0.0550 0.0300 ;
  LAYER VIA3 ;
    RECT -0.0250 -0.0250 0.0250 0.0250 ;
  LAYER M4 ;
    RECT -0.0300 -0.0550 0.0300 0.0550 ;
END VIA34SQ_C

VIA VIA34BAR_C
  RESISTANCE 1.6 ;
  LAYER M3 ;
    RECT -0.0550 -0.0550 0.0550 0.0550 ;
  LAYER VIA3 ;
    RECT -0.0250 -0.0500 0.0250 0.0500 ;
  LAYER M4 ;
    RECT -0.0300 -0.0800 0.0300 0.0800 ;
END VIA34BAR_C

VIA VIA34LG_C
  RESISTANCE 1.6 ;
  LAYER M3 ;
    RECT -0.0800 -0.0550 0.0800 0.0550 ;
  LAYER VIA3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M4 ;
    RECT -0.0800 -0.0550 0.0800 0.0550 ;
END VIA34LG_C

VIA VIA34SQ
  RESISTANCE 1.6 ;
  LAYER M3 ;
    RECT -0.0550 -0.0300 0.0550 0.0300 ;
  LAYER VIA3 ;
    RECT -0.0250 -0.0250 0.0250 0.0250 ;
  LAYER M4 ;
    RECT -0.0550 -0.0300 0.0550 0.0300 ;
END VIA34SQ

VIA VIA34BAR
  RESISTANCE 1.6 ;
  LAYER M3 ;
    RECT -0.0550 -0.0550 0.0550 0.0550 ;
  LAYER VIA3 ;
    RECT -0.0250 -0.0500 0.0250 0.0500 ;
  LAYER M4 ;
    RECT -0.0550 -0.0550 0.0550 0.0550 ;
END VIA34BAR

VIA VIA34LG
  RESISTANCE 1.6 ;
  LAYER M3 ;
    RECT -0.0800 -0.0550 0.0800 0.0550 ;
  LAYER VIA3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M4 ;
    RECT -0.0800 -0.0550 0.0800 0.0550 ;
END VIA34LG

VIA VIA45SQ_C
  DEFAULT 
  RESISTANCE 1.6 ;
  LAYER M4 ;
    RECT -0.0550 -0.0300 0.0550 0.0300 ;
  LAYER VIA4 ;
    RECT -0.0250 -0.0250 0.0250 0.0250 ;
  LAYER M5 ;
    RECT -0.0300 -0.0550 0.0300 0.0550 ;
END VIA45SQ_C

VIA VIA45BAR_C
  RESISTANCE 1.6 ;
  LAYER M4 ;
    RECT -0.0550 -0.0550 0.0550 0.0550 ;
  LAYER VIA4 ;
    RECT -0.0250 -0.0500 0.0250 0.0500 ;
  LAYER M5 ;
    RECT -0.0300 -0.0800 0.0300 0.0800 ;
END VIA45BAR_C

VIA VIA45LG_C
  RESISTANCE 1.6 ;
  LAYER M4 ;
    RECT -0.0800 -0.0550 0.0800 0.0550 ;
  LAYER VIA4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M5 ;
    RECT -0.0800 -0.0550 0.0800 0.0550 ;
END VIA45LG_C

VIA VIA45SQ
  RESISTANCE 1.6 ;
  LAYER M4 ;
    RECT -0.0550 -0.0300 0.0550 0.0300 ;
  LAYER VIA4 ;
    RECT -0.0250 -0.0250 0.0250 0.0250 ;
  LAYER M5 ;
    RECT -0.0550 -0.0300 0.0550 0.0300 ;
END VIA45SQ

VIA VIA45BAR
  RESISTANCE 1.6 ;
  LAYER M4 ;
    RECT -0.0550 -0.0550 0.0550 0.0550 ;
  LAYER VIA4 ;
    RECT -0.0250 -0.0500 0.0250 0.0500 ;
  LAYER M5 ;
    RECT -0.0550 -0.0550 0.0550 0.0550 ;
END VIA45BAR

VIA VIA45LG
  RESISTANCE 1.6 ;
  LAYER M4 ;
    RECT -0.0800 -0.0550 0.0800 0.0550 ;
  LAYER VIA4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M5 ;
    RECT -0.0800 -0.0550 0.0800 0.0550 ;
END VIA45LG

VIA VIA56SQ_C
  DEFAULT 
  RESISTANCE 1.6 ;
  LAYER M5 ;
    RECT -0.0550 -0.0300 0.0550 0.0300 ;
  LAYER VIA5 ;
    RECT -0.0250 -0.0250 0.0250 0.0250 ;
  LAYER M6 ;
    RECT -0.0300 -0.0550 0.0300 0.0550 ;
END VIA56SQ_C

VIA VIA56BAR_C
  RESISTANCE 1.6 ;
  LAYER M5 ;
    RECT -0.0550 -0.0550 0.0550 0.0550 ;
  LAYER VIA5 ;
    RECT -0.0250 -0.0500 0.0250 0.0500 ;
  LAYER M6 ;
    RECT -0.0300 -0.0800 0.0300 0.0800 ;
END VIA56BAR_C

VIA VIA56LG_C
  RESISTANCE 1.6 ;
  LAYER M5 ;
    RECT -0.0800 -0.0550 0.0800 0.0550 ;
  LAYER VIA5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M6 ;
    RECT -0.0800 -0.0550 0.0800 0.0550 ;
END VIA56LG_C

VIA VIA56SQ
  RESISTANCE 1.6 ;
  LAYER M5 ;
    RECT -0.0550 -0.0300 0.0550 0.0300 ;
  LAYER VIA5 ;
    RECT -0.0250 -0.0250 0.0250 0.0250 ;
  LAYER M6 ;
    RECT -0.0550 -0.0300 0.0550 0.0300 ;
END VIA56SQ

VIA VIA56BAR
  RESISTANCE 1.6 ;
  LAYER M5 ;
    RECT -0.0550 -0.0550 0.0550 0.0550 ;
  LAYER VIA5 ;
    RECT -0.0250 -0.0500 0.0250 0.0500 ;
  LAYER M6 ;
    RECT -0.0550 -0.0550 0.0550 0.0550 ;
END VIA56BAR

VIA VIA56LG
  RESISTANCE 1.6 ;
  LAYER M5 ;
    RECT -0.0800 -0.0550 0.0800 0.0550 ;
  LAYER VIA5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M6 ;
    RECT -0.0800 -0.0550 0.0800 0.0550 ;
END VIA56LG

VIA VIA67SQ_C
  DEFAULT 
  RESISTANCE 1.6 ;
  LAYER M6 ;
    RECT -0.0550 -0.0300 0.0550 0.0300 ;
  LAYER VIA6 ;
    RECT -0.0250 -0.0250 0.0250 0.0250 ;
  LAYER M7 ;
    RECT -0.0300 -0.0550 0.0300 0.0550 ;
END VIA67SQ_C

VIA VIA67BAR_C
  RESISTANCE 1.6 ;
  LAYER M6 ;
    RECT -0.0550 -0.0550 0.0550 0.0550 ;
  LAYER VIA6 ;
    RECT -0.0250 -0.0500 0.0250 0.0500 ;
  LAYER M7 ;
    RECT -0.0300 -0.0800 0.0300 0.0800 ;
END VIA67BAR_C

VIA VIA67LG_C
  RESISTANCE 1.6 ;
  LAYER M6 ;
    RECT -0.0800 -0.0550 0.0800 0.0550 ;
  LAYER VIA6 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M7 ;
    RECT -0.0800 -0.0550 0.0800 0.0550 ;
END VIA67LG_C

VIA VIA67SQ
  RESISTANCE 1.6 ;
  LAYER M6 ;
    RECT -0.0550 -0.0300 0.0550 0.0300 ;
  LAYER VIA6 ;
    RECT -0.0250 -0.0250 0.0250 0.0250 ;
  LAYER M7 ;
    RECT -0.0550 -0.0300 0.0550 0.0300 ;
END VIA67SQ

VIA VIA67BAR
  RESISTANCE 1.6 ;
  LAYER M6 ;
    RECT -0.0550 -0.0550 0.0550 0.0550 ;
  LAYER VIA6 ;
    RECT -0.0250 -0.0500 0.0250 0.0500 ;
  LAYER M7 ;
    RECT -0.0550 -0.0550 0.0550 0.0550 ;
END VIA67BAR

VIA VIA67LG
  RESISTANCE 1.6 ;
  LAYER M6 ;
    RECT -0.0800 -0.0550 0.0800 0.0550 ;
  LAYER VIA6 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M7 ;
    RECT -0.0800 -0.0550 0.0800 0.0550 ;
END VIA67LG

VIA VIA78SQ_C
  DEFAULT 
  RESISTANCE 1.6 ;
  LAYER M7 ;
    RECT -0.0550 -0.0300 0.0550 0.0300 ;
  LAYER VIA7 ;
    RECT -0.0250 -0.0250 0.0250 0.0250 ;
  LAYER M8 ;
    RECT -0.0300 -0.0550 0.0300 0.0550 ;
END VIA78SQ_C

VIA VIA78BAR_C
  RESISTANCE 1.6 ;
  LAYER M7 ;
    RECT -0.0550 -0.0550 0.0550 0.0550 ;
  LAYER VIA7 ;
    RECT -0.0250 -0.0500 0.0250 0.0500 ;
  LAYER M8 ;
    RECT -0.0300 -0.0800 0.0300 0.0800 ;
END VIA78BAR_C

VIA VIA78LG_C
  RESISTANCE 1.6 ;
  LAYER M7 ;
    RECT -0.0800 -0.0550 0.0800 0.0550 ;
  LAYER VIA7 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M8 ;
    RECT -0.0800 -0.0550 0.0800 0.0550 ;
END VIA78LG_C

VIA VIA78SQ
  RESISTANCE 1.6 ;
  LAYER M7 ;
    RECT -0.0550 -0.0300 0.0550 0.0300 ;
  LAYER VIA7 ;
    RECT -0.0250 -0.0250 0.0250 0.0250 ;
  LAYER M8 ;
    RECT -0.0550 -0.0300 0.0550 0.0300 ;
END VIA78SQ

VIA VIA78BAR
  RESISTANCE 1.6 ;
  LAYER M7 ;
    RECT -0.0550 -0.0550 0.0550 0.0550 ;
  LAYER VIA7 ;
    RECT -0.0250 -0.0500 0.0250 0.0500 ;
  LAYER M8 ;
    RECT -0.0550 -0.0550 0.0550 0.0550 ;
END VIA78BAR

VIA VIA78LG
  RESISTANCE 1.6 ;
  LAYER M7 ;
    RECT -0.0800 -0.0550 0.0800 0.0550 ;
  LAYER VIA7 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
  LAYER M8 ;
    RECT -0.0800 -0.0550 0.0800 0.0550 ;
END VIA78LG

VIA VIA89_C
  DEFAULT 
  RESISTANCE 1.6 ;
  LAYER M8 ;
    RECT -0.0950 -0.0800 0.0950 0.0800 ;
  LAYER VIA8 ;
    RECT -0.0650 -0.0650 0.0650 0.0650 ;
  LAYER M9 ;
    RECT -0.0800 -0.0950 0.0800 0.0950 ;
END VIA89_C

VIA VIA89
  DEFAULT 
  RESISTANCE 1.6 ;
  LAYER M8 ;
    RECT -0.0950 -0.0800 0.0950 0.0800 ;
  LAYER VIA8 ;
    RECT -0.0650 -0.0650 0.0650 0.0650 ;
  LAYER M9 ;
    RECT -0.0950 -0.0800 0.0950 0.0800 ;
END VIA89

VIA VIA9RDL
  DEFAULT 
  RESISTANCE 1.6 ;
  LAYER M9 ;
    RECT -1.5000 -1.5000 1.5000 1.5000 ;
  LAYER VIARDL ;
    RECT -1.0000 -1.0000 1.0000 1.0000 ;
  LAYER MRDL ;
    RECT -1.5000 -1.5000 1.5000 1.5000 ;
END VIA9RDL

VIARULE VIA12SQ_C GENERATE
  LAYER M1 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M2 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER VIA1 ;
    RECT -0.0250 -0.0250 0.0250 0.0250 ;
    SPACING 0.12 BY 0.12 ;
    RESISTANCE 1.6 ;
END VIA12SQ_C

VIARULE VIA12BAR_C GENERATE
  LAYER M1 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M2 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER VIA1 ;
    RECT -0.0250 -0.0500 0.0250 0.0500 ;
    SPACING 0.135 BY 0.185 ;
    RESISTANCE 1.6 ;
END VIA12BAR_C

VIARULE VIA12LG_C GENERATE
  LAYER M1 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
  LAYER M2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.005 ;
  LAYER VIA1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.185 BY 0.185 ;
    RESISTANCE 1.6 ;
END VIA12LG_C

VIARULE VIA12SQ GENERATE
  LAYER M1 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
  LAYER M2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.005 ;
  LAYER VIA1 ;
    RECT -0.0250 -0.0250 0.0250 0.0250 ;
    SPACING 0.12 BY 0.12 ;
    RESISTANCE 1.6 ;
END VIA12SQ

VIARULE VIA12BAR GENERATE
  LAYER M1 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
  LAYER M2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.005 ;
  LAYER VIA1 ;
    RECT -0.0250 -0.0500 0.0250 0.0500 ;
    SPACING 0.135 BY 0.185 ;
    RESISTANCE 1.6 ;
END VIA12BAR

VIARULE VIA12LG GENERATE
  LAYER M1 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
  LAYER M2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.005 ;
  LAYER VIA1 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.185 BY 0.185 ;
    RESISTANCE 1.6 ;
END VIA12LG

VIARULE VIA23SQ_C GENERATE
  LAYER M2 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M3 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER VIA2 ;
    RECT -0.0250 -0.0250 0.0250 0.0250 ;
    SPACING 0.12 BY 0.12 ;
    RESISTANCE 1.6 ;
END VIA23SQ_C

VIARULE VIA23BAR_C GENERATE
  LAYER M2 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M3 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER VIA2 ;
    RECT -0.0250 -0.0500 0.0250 0.0500 ;
    SPACING 0.135 BY 0.185 ;
    RESISTANCE 1.6 ;
END VIA23BAR_C

VIARULE VIA23LG_C GENERATE
  LAYER M2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.005 ;
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
  LAYER VIA2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.185 BY 0.185 ;
    RESISTANCE 1.6 ;
END VIA23LG_C

VIARULE VIA23SQ GENERATE
  LAYER M2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.005 ;
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
  LAYER VIA2 ;
    RECT -0.0250 -0.0250 0.0250 0.0250 ;
    SPACING 0.12 BY 0.12 ;
    RESISTANCE 1.6 ;
END VIA23SQ

VIARULE VIA23BAR GENERATE
  LAYER M2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.005 ;
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
  LAYER VIA2 ;
    RECT -0.0250 -0.0500 0.0250 0.0500 ;
    SPACING 0.135 BY 0.185 ;
    RESISTANCE 1.6 ;
END VIA23BAR

VIARULE VIA23LG GENERATE
  LAYER M2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.005 ;
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
  LAYER VIA2 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.185 BY 0.185 ;
    RESISTANCE 1.6 ;
END VIA23LG

VIARULE VIA34SQ_C GENERATE
  LAYER M3 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M4 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER VIA3 ;
    RECT -0.0250 -0.0250 0.0250 0.0250 ;
    SPACING 0.12 BY 0.12 ;
    RESISTANCE 1.6 ;
END VIA34SQ_C

VIARULE VIA34BAR_C GENERATE
  LAYER M3 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M4 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER VIA3 ;
    RECT -0.0250 -0.0500 0.0250 0.0500 ;
    SPACING 0.135 BY 0.185 ;
    RESISTANCE 1.6 ;
END VIA34BAR_C

VIARULE VIA34LG_C GENERATE
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
  LAYER M4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.005 ;
  LAYER VIA3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.185 BY 0.185 ;
    RESISTANCE 1.6 ;
END VIA34LG_C

VIARULE VIA34SQ GENERATE
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
  LAYER M4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.005 ;
  LAYER VIA3 ;
    RECT -0.0250 -0.0250 0.0250 0.0250 ;
    SPACING 0.12 BY 0.12 ;
    RESISTANCE 1.6 ;
END VIA34SQ

VIARULE VIA34BAR GENERATE
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
  LAYER M4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.005 ;
  LAYER VIA3 ;
    RECT -0.0250 -0.0500 0.0250 0.0500 ;
    SPACING 0.135 BY 0.185 ;
    RESISTANCE 1.6 ;
END VIA34BAR

VIARULE VIA34LG GENERATE
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
  LAYER M4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.005 ;
  LAYER VIA3 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.185 BY 0.185 ;
    RESISTANCE 1.6 ;
END VIA34LG

VIARULE VIA45SQ_C GENERATE
  LAYER M4 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M5 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER VIA4 ;
    RECT -0.0250 -0.0250 0.0250 0.0250 ;
    SPACING 0.12 BY 0.12 ;
    RESISTANCE 1.6 ;
END VIA45SQ_C

VIARULE VIA45BAR_C GENERATE
  LAYER M4 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M5 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER VIA4 ;
    RECT -0.0250 -0.0500 0.0250 0.0500 ;
    SPACING 0.135 BY 0.185 ;
    RESISTANCE 1.6 ;
END VIA45BAR_C

VIARULE VIA45LG_C GENERATE
  LAYER M4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.005 ;
  LAYER M5 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
  LAYER VIA4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.185 BY 0.185 ;
    RESISTANCE 1.6 ;
END VIA45LG_C

VIARULE VIA45SQ GENERATE
  LAYER M4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.005 ;
  LAYER M5 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
  LAYER VIA4 ;
    RECT -0.0250 -0.0250 0.0250 0.0250 ;
    SPACING 0.12 BY 0.12 ;
    RESISTANCE 1.6 ;
END VIA45SQ

VIARULE VIA45BAR GENERATE
  LAYER M4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.005 ;
  LAYER M5 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
  LAYER VIA4 ;
    RECT -0.0250 -0.0500 0.0250 0.0500 ;
    SPACING 0.135 BY 0.185 ;
    RESISTANCE 1.6 ;
END VIA45BAR

VIARULE VIA45LG GENERATE
  LAYER M4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.005 ;
  LAYER M5 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
  LAYER VIA4 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.185 BY 0.185 ;
    RESISTANCE 1.6 ;
END VIA45LG

VIARULE VIA56SQ_C GENERATE
  LAYER M5 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M6 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER VIA5 ;
    RECT -0.0250 -0.0250 0.0250 0.0250 ;
    SPACING 0.12 BY 0.12 ;
    RESISTANCE 1.6 ;
END VIA56SQ_C

VIARULE VIA56BAR_C GENERATE
  LAYER M5 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M6 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER VIA5 ;
    RECT -0.0250 -0.0500 0.0250 0.0500 ;
    SPACING 0.135 BY 0.185 ;
    RESISTANCE 1.6 ;
END VIA56BAR_C

VIARULE VIA56LG_C GENERATE
  LAYER M5 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
  LAYER M6 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.005 ;
  LAYER VIA5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.185 BY 0.185 ;
    RESISTANCE 1.6 ;
END VIA56LG_C

VIARULE VIA56SQ GENERATE
  LAYER M5 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
  LAYER M6 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.005 ;
  LAYER VIA5 ;
    RECT -0.0250 -0.0250 0.0250 0.0250 ;
    SPACING 0.12 BY 0.12 ;
    RESISTANCE 1.6 ;
END VIA56SQ

VIARULE VIA56BAR GENERATE
  LAYER M5 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
  LAYER M6 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.005 ;
  LAYER VIA5 ;
    RECT -0.0250 -0.0500 0.0250 0.0500 ;
    SPACING 0.135 BY 0.185 ;
    RESISTANCE 1.6 ;
END VIA56BAR

VIARULE VIA56LG GENERATE
  LAYER M5 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
  LAYER M6 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.005 ;
  LAYER VIA5 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.185 BY 0.185 ;
    RESISTANCE 1.6 ;
END VIA56LG

VIARULE VIA67SQ_C GENERATE
  LAYER M6 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M7 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER VIA6 ;
    RECT -0.0250 -0.0250 0.0250 0.0250 ;
    SPACING 0.12 BY 0.12 ;
    RESISTANCE 1.6 ;
END VIA67SQ_C

VIARULE VIA67BAR_C GENERATE
  LAYER M6 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M7 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER VIA6 ;
    RECT -0.0250 -0.0500 0.0250 0.0500 ;
    SPACING 0.135 BY 0.185 ;
    RESISTANCE 1.6 ;
END VIA67BAR_C

VIARULE VIA67LG_C GENERATE
  LAYER M6 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.005 ;
  LAYER M7 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
  LAYER VIA6 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.185 BY 0.185 ;
    RESISTANCE 1.6 ;
END VIA67LG_C

VIARULE VIA67SQ GENERATE
  LAYER M6 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.005 ;
  LAYER M7 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
  LAYER VIA6 ;
    RECT -0.0250 -0.0250 0.0250 0.0250 ;
    SPACING 0.12 BY 0.12 ;
    RESISTANCE 1.6 ;
END VIA67SQ

VIARULE VIA67BAR GENERATE
  LAYER M6 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.005 ;
  LAYER M7 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
  LAYER VIA6 ;
    RECT -0.0250 -0.0500 0.0250 0.0500 ;
    SPACING 0.135 BY 0.185 ;
    RESISTANCE 1.6 ;
END VIA67BAR

VIARULE VIA67LG GENERATE
  LAYER M6 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.005 ;
  LAYER M7 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
  LAYER VIA6 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.185 BY 0.185 ;
    RESISTANCE 1.6 ;
END VIA67LG

VIARULE VIA78SQ_C GENERATE
  LAYER M7 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M8 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER VIA7 ;
    RECT -0.0250 -0.0250 0.0250 0.0250 ;
    SPACING 0.12 BY 0.12 ;
    RESISTANCE 1.6 ;
END VIA78SQ_C

VIARULE VIA78BAR_C GENERATE
  LAYER M7 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M8 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER VIA7 ;
    RECT -0.0250 -0.0500 0.0250 0.0500 ;
    SPACING 0.135 BY 0.185 ;
    RESISTANCE 1.6 ;
END VIA78BAR_C

VIARULE VIA78LG_C GENERATE
  LAYER M7 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
  LAYER M8 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.005 ;
  LAYER VIA7 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.185 BY 0.185 ;
    RESISTANCE 1.6 ;
END VIA78LG_C

VIARULE VIA78SQ GENERATE
  LAYER M7 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
  LAYER M8 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.005 ;
  LAYER VIA7 ;
    RECT -0.0250 -0.0250 0.0250 0.0250 ;
    SPACING 0.12 BY 0.12 ;
    RESISTANCE 1.6 ;
END VIA78SQ

VIARULE VIA78BAR GENERATE
  LAYER M7 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
  LAYER M8 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.005 ;
  LAYER VIA7 ;
    RECT -0.0250 -0.0500 0.0250 0.0500 ;
    SPACING 0.135 BY 0.185 ;
    RESISTANCE 1.6 ;
END VIA78BAR

VIARULE VIA78LG GENERATE
  LAYER M7 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
  LAYER M8 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.005 ;
  LAYER VIA7 ;
    RECT -0.0500 -0.0500 0.0500 0.0500 ;
    SPACING 0.185 BY 0.185 ;
    RESISTANCE 1.6 ;
END VIA78LG

VIARULE VIA89_C GENERATE
  LAYER M8 ;
    ENCLOSURE 0.03 0.015 ;
  LAYER M9 ;
    ENCLOSURE 0.015 0.03 ;
  LAYER VIA8 ;
    RECT -0.0650 -0.0650 0.0650 0.0650 ;
    SPACING 0.25 BY 0.25 ;
    RESISTANCE 1.6 ;
END VIA89_C

VIARULE VIA89 GENERATE
  LAYER M8 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.015 ;
  LAYER M9 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
  LAYER VIA8 ;
    RECT -0.0650 -0.0650 0.0650 0.0650 ;
    SPACING 0.25 BY 0.25 ;
    RESISTANCE 1.6 ;
END VIA89

VIARULE VIA9RDL GENERATE
  LAYER M9 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.5 ;
  LAYER MRDL ;
    DIRECTION VERTICAL ;
    OVERHANG 0.5 ;
  LAYER VIARDL ;
    RECT -1.0000 -1.0000 1.0000 1.0000 ;
    SPACING 4 BY 4 ;
    RESISTANCE 1.6 ;
END VIA9RDL


SITE ioSiteNS
  CLASS PAD ;
  SYMMETRY R90 ;
  SIZE 0.1 BY 300 ;
END ioSiteNS

SITE ioSiteEW
  CLASS PAD ;
  SYMMETRY R90 ;
  SIZE 300 BY 0.1 ;
END ioSiteEW

SITE cornerSite
  CLASS PAD ;
  SYMMETRY R90 ;
  SIZE 300 BY 300 ;
END cornerSite

SITE fillSite 
  CLASS PAD ;
  SYMMETRY R90 ;
  SIZE 300 BY 0.1 ;
END fillSite

SITE unit
  CLASS CORE ;
  SYMMETRY X Y ;
  SIZE 0.152 BY 1.672 ;
END unit

  
END LIBRARY
