#######################################################################
####                                                               ####
####  The data contained in the file is created for educational    #### 
####  and training purposes only and are not recommended           ####
####  for fabrication                                              ####
####                                                               ####
#######################################################################
####                                                               ####
####  Copyright (C) 2013 Synopsys, Inc.                            ####
####                                                               ####
#######################################################################
####                                                               ####
####  The 32/28nm Generic Library ("Library") is unsupported       ####    
####  Confidential Information of Synopsys, Inc. ("Synopsys")      ####    
####  provided to you as Documentation under the terms of the      ####    
####  End User Software License Agreement between you or your      ####    
####  employer and Synopsys ("License Agreement") and you agree    ####    
####  not to distribute or disclose the Library without the        ####    
####  prior written consent of Synopsys. The Library IS NOT an     ####    
####  item of Licensed Software or Licensed Product under the      ####    
####  License Agreement.  Synopsys and/or its licensors own        ####    
####  and shall retain all right, title and interest in and        ####    
####  to the Library and all modifications thereto, including      ####    
####  all intellectual property rights embodied therein. All       ####    
####  rights in and to any Library modifications you make are      ####    
####  hereby assigned to Synopsys. If you do not agree with        ####    
####  this notice, including the disclaimer below, then you        ####    
####  are not authorized to use the Library.                       ####    
####                                                               ####  
####                                                               ####      
####  THIS LIBRARY IS BEING DISTRIBUTED BY SYNOPSYS SOLELY ON AN   ####
####  "AS IS" BASIS, WITH NO INTELLECUTAL PROPERTY                 ####
####  INDEMNIFICATION AND NO SUPPORT. ANY EXPRESS OR IMPLIED       ####
####  WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED       ####
####  WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR   ####
####  PURPOSE ARE HEREBY DISCLAIMED. IN NO EVENT SHALL SYNOPSYS    ####
####  BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL,     ####
####  EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT      ####
####  LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;     ####
####  LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)     ####
####  HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN    ####
####  CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE    ####
####  OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS      ####
####  DOCUMENTATION, EVEN IF ADVISED OF THE POSSIBILITY OF         ####
####  SUCH DAMAGE.                                                 #### 
####                                                               ####  
#######################################################################

# 
# LEF OUT 
# User Name : edbab 
# Date : Mon Dec 24 17:39:53 2012
# 
VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;

MACRO TNBUFFX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.128 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3240 1.3730 0.7360 1.4230 ;
        RECT 0.5530 1.4230 0.6630 1.5750 ;
    END
    ANTENNAGATEAREA 0.0264 ;
  END EN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.1280 1.7020 ;
        RECT 1.6470 1.2720 1.6970 1.6420 ;
        RECT 0.2240 1.2060 0.2740 1.6420 ;
        RECT 0.8100 1.1100 0.8600 1.6420 ;
        RECT 0.2240 1.1560 0.3290 1.2060 ;
        RECT 0.7350 1.0600 0.9370 1.1100 ;
        RECT 0.2790 0.7310 0.3290 1.1560 ;
        RECT 0.7350 0.8140 0.7850 1.0600 ;
        RECT 0.8870 0.8140 0.9370 1.0600 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.1280 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.5420 ;
        RECT 1.6470 0.0300 1.6970 0.1880 ;
        RECT 1.0390 0.1880 1.6970 0.2380 ;
        RECT 1.0390 0.2380 1.0890 0.5520 ;
        RECT 1.1920 0.2380 1.2420 0.5520 ;
        RECT 1.6470 0.2380 1.6970 0.3680 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8540 0.4870 1.9040 0.6780 ;
        RECT 1.8540 0.6780 2.0510 0.8150 ;
        RECT 1.4950 0.4370 1.9040 0.4870 ;
        RECT 1.8540 0.8150 1.9040 1.0840 ;
        RECT 1.7990 0.1110 1.8490 0.4370 ;
        RECT 1.4950 0.2880 1.5450 0.4370 ;
        RECT 1.4950 1.0840 1.9040 1.1340 ;
        RECT 1.7990 1.1340 1.8490 1.4720 ;
        RECT 1.4950 1.1340 1.5450 1.4720 ;
    END
    ANTENNADIFFAREA 0.2222 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9320 1.4030 1.1190 1.4530 ;
        RECT 1.0090 1.3130 1.1190 1.4030 ;
    END
    ANTENNAGATEAREA 0.0243 ;
  END A
  OBS
    LAYER NWELL ;
      RECT -0.1120 0.6790 2.2400 1.7730 ;
    LAYER M1 ;
      RECT 1.4570 0.5570 1.8040 0.5870 ;
      RECT 1.4580 0.5370 1.8040 0.5570 ;
      RECT 0.8120 0.5510 0.8620 0.6020 ;
      RECT 0.7350 0.5010 0.9370 0.5510 ;
      RECT 0.8870 0.3430 0.9370 0.5010 ;
      RECT 0.7350 0.3430 0.7850 0.5010 ;
      RECT 1.3430 0.6520 1.3930 0.9340 ;
      RECT 1.3430 0.3480 1.3930 0.6020 ;
      RECT 1.4570 0.5870 1.5070 0.6020 ;
      RECT 0.8120 0.6020 1.5070 0.6520 ;
      RECT 1.5400 0.7450 1.8040 0.7950 ;
      RECT 0.5830 0.3480 0.6330 0.7140 ;
      RECT 0.5830 0.7640 0.6330 1.0180 ;
      RECT 1.0390 0.7640 1.0890 1.2020 ;
      RECT 1.1920 0.7640 1.2420 0.9840 ;
      RECT 1.1920 0.7130 1.2420 0.7140 ;
      RECT 0.5830 0.7140 1.2420 0.7640 ;
      RECT 1.5710 0.7950 1.6210 0.9840 ;
      RECT 1.1920 0.9840 1.6210 1.0340 ;
      RECT 0.4310 0.0880 1.3480 0.1380 ;
      RECT 0.4310 0.1380 0.4810 1.1190 ;
    LAYER PO ;
      RECT 1.5810 0.0660 1.6110 0.6150 ;
      RECT 1.5810 0.7170 1.6110 1.6060 ;
      RECT 1.7330 0.0660 1.7630 0.6150 ;
      RECT 1.7330 0.7170 1.7630 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
  END
END TNBUFFX2_LVT

MACRO TNBUFFX32_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.488 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0970 0.5530 0.2070 0.6020 ;
        RECT 0.0970 0.6020 0.4360 0.6520 ;
        RECT 0.0970 0.6520 0.2070 0.6630 ;
    END
    ANTENNAGATEAREA 0.0264 ;
  END A

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0990 0.6600 1.3330 0.7100 ;
        RECT 1.1610 0.7100 1.2710 0.8150 ;
    END
    ANTENNAGATEAREA 0.0732 ;
  END EN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 10.4880 1.7020 ;
        RECT 1.6020 1.4690 1.6520 1.6420 ;
        RECT 1.1910 1.4190 1.6970 1.4690 ;
        RECT 5.4470 1.2750 5.4970 1.6420 ;
        RECT 5.7510 1.2720 5.8010 1.6420 ;
        RECT 6.0550 1.2720 6.1050 1.6420 ;
        RECT 6.3590 1.2720 6.4090 1.6420 ;
        RECT 6.6630 1.2720 6.7130 1.6420 ;
        RECT 6.9670 1.2720 7.0170 1.6420 ;
        RECT 7.2710 1.2720 7.3210 1.6420 ;
        RECT 7.5750 1.2720 7.6250 1.6420 ;
        RECT 7.8790 1.2750 7.9290 1.6420 ;
        RECT 8.1830 1.2720 8.2330 1.6420 ;
        RECT 8.4870 1.2720 8.5370 1.6420 ;
        RECT 8.7910 1.2720 8.8410 1.6420 ;
        RECT 9.0950 1.2720 9.1450 1.6420 ;
        RECT 9.3990 1.2720 9.4490 1.6420 ;
        RECT 9.7030 1.2720 9.7530 1.6420 ;
        RECT 10.0070 1.2720 10.0570 1.6420 ;
        RECT 4.1340 1.3130 4.1840 1.6420 ;
        RECT 0.7350 0.9350 0.7850 1.6420 ;
        RECT 0.2790 0.7460 0.3290 1.6420 ;
        RECT 3.9270 1.3130 3.9770 1.4940 ;
        RECT 3.6230 1.3130 3.6730 1.4940 ;
        RECT 3.3190 1.3130 3.3690 1.4940 ;
        RECT 1.1910 1.2950 1.2410 1.4190 ;
        RECT 1.6470 1.2950 1.6970 1.4190 ;
        RECT 2.1030 1.2630 4.1840 1.3130 ;
        RECT 2.4070 0.9380 2.4570 1.2630 ;
        RECT 2.7110 0.9380 2.7610 1.2630 ;
        RECT 2.1030 0.9380 2.1530 1.2630 ;
        RECT 3.9270 0.8600 3.9770 1.2630 ;
        RECT 3.6230 0.8600 3.6730 1.2630 ;
        RECT 3.3190 0.8600 3.3690 1.2630 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 10.4880 0.0300 ;
        RECT 5.7510 0.0300 5.8010 0.3380 ;
        RECT 7.5750 0.0300 7.6250 0.3380 ;
        RECT 7.2710 0.0300 7.3210 0.3380 ;
        RECT 6.9670 0.0300 7.0170 0.3380 ;
        RECT 6.6630 0.0300 6.7130 0.3380 ;
        RECT 1.1910 0.0300 1.2410 0.3800 ;
        RECT 6.3590 0.0300 6.4090 0.3380 ;
        RECT 6.0550 0.0300 6.1050 0.3380 ;
        RECT 0.2790 0.0300 0.3290 0.4720 ;
        RECT 0.7350 0.0300 0.7850 0.3270 ;
        RECT 1.6470 0.0300 1.6970 0.2230 ;
        RECT 7.8790 0.0300 7.9290 0.3380 ;
        RECT 8.1830 0.0300 8.2330 0.3380 ;
        RECT 10.0070 0.0300 10.0570 0.3380 ;
        RECT 9.7030 0.0300 9.7530 0.3380 ;
        RECT 9.3990 0.0300 9.4490 0.3380 ;
        RECT 9.0950 0.0300 9.1450 0.3380 ;
        RECT 8.7910 0.0300 8.8410 0.3380 ;
        RECT 8.4870 0.0300 8.5370 0.3380 ;
        RECT 5.4470 0.0300 5.4970 0.2050 ;
        RECT 3.1670 0.2050 5.4970 0.2550 ;
        RECT 3.1670 0.2550 3.2170 0.3950 ;
        RECT 4.9920 0.2550 5.0420 0.4450 ;
        RECT 3.4710 0.2550 3.5210 0.3950 ;
        RECT 3.7750 0.2550 3.8250 0.3950 ;
        RECT 4.0790 0.2550 4.1290 0.3950 ;
        RECT 4.3840 0.2550 4.4340 0.4450 ;
        RECT 4.6880 0.2550 4.7380 0.4450 ;
        RECT 5.4470 0.2550 5.4970 0.3380 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.2470 1.1340 9.2970 1.5090 ;
        RECT 9.5510 1.1340 9.6010 1.5090 ;
        RECT 9.8550 1.1340 9.9050 1.5090 ;
        RECT 10.1590 1.1340 10.2090 1.4720 ;
        RECT 8.0310 1.1340 8.0810 1.5090 ;
        RECT 8.3350 1.1340 8.3850 1.5090 ;
        RECT 8.6390 1.1340 8.6890 1.5090 ;
        RECT 8.9430 1.1340 8.9930 1.5090 ;
        RECT 6.8150 1.1340 6.8650 1.5090 ;
        RECT 7.1190 1.1340 7.1690 1.5090 ;
        RECT 7.4230 1.1340 7.4730 1.5090 ;
        RECT 7.7270 1.1340 7.7770 1.5090 ;
        RECT 5.2950 1.1340 5.3450 1.5090 ;
        RECT 5.5990 1.1340 5.6490 1.5090 ;
        RECT 5.9030 1.1340 5.9530 1.5090 ;
        RECT 6.2070 1.1340 6.2570 1.5090 ;
        RECT 6.5110 1.1340 6.5610 1.5090 ;
        RECT 5.2950 1.0840 10.2640 1.1340 ;
        RECT 10.2140 0.9670 10.2640 1.0840 ;
        RECT 9.2470 0.8450 9.2970 1.0840 ;
        RECT 9.5510 0.8450 9.6010 1.0840 ;
        RECT 9.8550 0.8450 9.9050 1.0840 ;
        RECT 10.2140 0.8570 10.3910 0.9670 ;
        RECT 8.0310 0.8450 8.0810 1.0840 ;
        RECT 8.3350 0.8450 8.3850 1.0840 ;
        RECT 8.6390 0.8450 8.6890 1.0840 ;
        RECT 8.9430 0.8450 8.9930 1.0840 ;
        RECT 7.4230 0.8450 7.4730 1.0840 ;
        RECT 6.8150 0.8450 6.8650 1.0840 ;
        RECT 7.1190 0.8450 7.1690 1.0840 ;
        RECT 7.7270 0.8450 7.7770 1.0840 ;
        RECT 5.5990 0.8450 5.6490 1.0840 ;
        RECT 5.9030 0.8450 5.9530 1.0840 ;
        RECT 6.2070 0.8450 6.2570 1.0840 ;
        RECT 6.5110 0.8450 6.5610 1.0840 ;
        RECT 5.2950 0.3880 10.2640 0.4380 ;
        RECT 8.0310 0.1420 8.0810 0.3880 ;
        RECT 8.3350 0.1420 8.3850 0.3880 ;
        RECT 8.6390 0.1420 8.6890 0.3880 ;
        RECT 8.9430 0.1420 8.9930 0.3880 ;
        RECT 10.2140 0.4380 10.2640 0.8570 ;
        RECT 9.2470 0.1420 9.2970 0.3880 ;
        RECT 9.5510 0.1420 9.6010 0.3880 ;
        RECT 9.8550 0.1420 9.9050 0.3880 ;
        RECT 10.1590 0.1420 10.2090 0.3880 ;
        RECT 6.8150 0.1420 6.8650 0.3880 ;
        RECT 7.1190 0.1420 7.1690 0.3880 ;
        RECT 7.4230 0.1420 7.4730 0.3880 ;
        RECT 7.7270 0.1420 7.7770 0.3880 ;
        RECT 5.5990 0.1420 5.6490 0.3880 ;
        RECT 5.9030 0.1420 5.9530 0.3880 ;
        RECT 6.2070 0.1420 6.2570 0.3880 ;
        RECT 6.5110 0.1420 6.5610 0.3880 ;
        RECT 5.2950 0.3560 5.3450 0.3880 ;
    END
    ANTENNADIFFAREA 2.2151 ;
  END Y
  OBS
    LAYER PO ;
      RECT 8.4210 0.7170 8.4510 1.6060 ;
      RECT 10.0930 0.0660 10.1230 0.6170 ;
      RECT 9.7890 0.0660 9.8190 0.6170 ;
      RECT 9.6370 0.0660 9.6670 0.6170 ;
      RECT 9.9410 0.0660 9.9710 0.6170 ;
      RECT 9.4850 0.0660 9.5150 0.6170 ;
      RECT 9.3330 0.0660 9.3630 0.6170 ;
      RECT 9.1810 0.0660 9.2110 0.6170 ;
      RECT 9.0290 0.0660 9.0590 0.6170 ;
      RECT 8.5730 0.0660 8.6030 0.6170 ;
      RECT 8.8770 0.0660 8.9070 0.6170 ;
      RECT 8.7250 0.0660 8.7550 0.6170 ;
      RECT 8.4210 0.0660 8.4510 0.6170 ;
      RECT 7.6610 0.0660 7.6910 0.6170 ;
      RECT 7.6610 0.7170 7.6910 1.6060 ;
      RECT 7.3570 0.0660 7.3870 0.6170 ;
      RECT 7.3570 0.7170 7.3870 1.6060 ;
      RECT 7.2050 0.0660 7.2350 0.6170 ;
      RECT 7.2050 0.7170 7.2350 1.6060 ;
      RECT 7.5090 0.0660 7.5390 0.6170 ;
      RECT 7.5090 0.7170 7.5390 1.6060 ;
      RECT 7.0530 0.0660 7.0830 0.6170 ;
      RECT 7.0530 0.7170 7.0830 1.6060 ;
      RECT 6.9010 0.0660 6.9310 0.6170 ;
      RECT 6.9010 0.7170 6.9310 1.6060 ;
      RECT 6.7490 0.0660 6.7790 0.6170 ;
      RECT 6.7490 0.7170 6.7790 1.6060 ;
      RECT 6.5970 0.0660 6.6270 0.6170 ;
      RECT 6.5970 0.7170 6.6270 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 6.1410 0.0660 6.1710 0.6170 ;
      RECT 6.1410 0.7170 6.1710 1.6060 ;
      RECT 6.4450 0.0660 6.4750 0.6170 ;
      RECT 6.4450 0.7170 6.4750 1.6060 ;
      RECT 6.2930 0.0660 6.3230 0.6170 ;
      RECT 6.2930 0.7170 6.3230 1.6060 ;
      RECT 5.9890 0.0660 6.0190 0.6170 ;
      RECT 5.9890 0.7170 6.0190 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 5.5330 0.7170 5.5630 1.6060 ;
      RECT 5.6850 0.7170 5.7150 1.6060 ;
      RECT 5.8370 0.7170 5.8670 1.6060 ;
      RECT 5.3810 0.7170 5.4110 1.6060 ;
      RECT 5.3810 0.0660 5.4110 0.6170 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 5.8370 0.0660 5.8670 0.6170 ;
      RECT 5.6850 0.0660 5.7150 0.6170 ;
      RECT 5.5330 0.0660 5.5630 0.6170 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 3.7090 0.0660 3.7390 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 10.3970 0.0660 10.4270 1.6060 ;
      RECT 10.2450 0.0660 10.2750 1.6060 ;
      RECT 7.9650 0.7170 7.9950 1.6060 ;
      RECT 8.1170 0.7170 8.1470 1.6060 ;
      RECT 8.2690 0.7170 8.2990 1.6060 ;
      RECT 7.8130 0.7170 7.8430 1.6060 ;
      RECT 7.8130 0.0660 7.8430 0.6170 ;
      RECT 8.2690 0.0660 8.2990 0.6170 ;
      RECT 8.1170 0.0660 8.1470 0.6170 ;
      RECT 7.9650 0.0660 7.9950 0.6170 ;
      RECT 10.0930 0.7170 10.1230 1.6060 ;
      RECT 9.7890 0.7170 9.8190 1.6060 ;
      RECT 9.6370 0.7170 9.6670 1.6060 ;
      RECT 9.9410 0.7170 9.9710 1.6060 ;
      RECT 9.4850 0.7170 9.5150 1.6060 ;
      RECT 9.3330 0.7170 9.3630 1.6060 ;
      RECT 9.1810 0.7170 9.2110 1.6060 ;
      RECT 9.0290 0.7170 9.0590 1.6060 ;
      RECT 8.5730 0.7170 8.6030 1.6060 ;
      RECT 8.8770 0.7170 8.9070 1.6060 ;
      RECT 8.7250 0.7170 8.7550 1.6060 ;
    LAYER NWELL ;
      RECT -0.1120 0.6790 10.6000 1.7730 ;
    LAYER M1 ;
      RECT 5.3400 0.7450 10.1640 0.7950 ;
      RECT 1.9510 0.8100 2.0010 1.3130 ;
      RECT 1.9510 0.2620 2.0010 0.7600 ;
      RECT 2.2550 0.2620 2.3050 0.4460 ;
      RECT 2.2550 0.8100 2.3050 1.2130 ;
      RECT 2.5590 0.2620 2.6090 0.4460 ;
      RECT 2.5590 0.8100 2.6090 1.2130 ;
      RECT 1.9510 0.2120 2.9130 0.2620 ;
      RECT 2.8630 0.2620 2.9130 0.4460 ;
      RECT 2.8630 0.8100 2.9130 1.2130 ;
      RECT 3.1670 0.8100 3.2170 1.2130 ;
      RECT 3.4710 0.8100 3.5210 1.2120 ;
      RECT 3.7750 0.8100 3.8250 1.2120 ;
      RECT 4.0790 0.8100 4.1290 1.1520 ;
      RECT 1.9500 0.7600 4.1290 0.8100 ;
      RECT 4.3840 0.8530 4.4340 1.1520 ;
      RECT 4.6880 0.8530 4.7380 1.1520 ;
      RECT 4.0790 1.1520 5.0420 1.2020 ;
      RECT 4.9920 1.0340 5.0420 1.1520 ;
      RECT 4.9920 0.8530 5.0420 0.9840 ;
      RECT 5.3400 0.7950 5.3900 0.9840 ;
      RECT 4.9920 0.9840 5.3900 1.0340 ;
      RECT 1.8490 1.3900 2.8680 1.4400 ;
      RECT 1.4950 0.8330 1.5450 0.9870 ;
      RECT 1.8490 0.8330 1.8990 1.3900 ;
      RECT 1.4950 0.7830 1.8990 0.8330 ;
      RECT 1.8490 0.4570 1.8990 0.7830 ;
      RECT 1.4640 0.4070 1.8990 0.4570 ;
      RECT 1.8330 0.1000 5.1480 0.1500 ;
      RECT 1.0390 0.1920 1.0890 0.5000 ;
      RECT 1.0390 0.9150 1.0890 1.1450 ;
      RECT 1.3430 0.3570 1.3930 0.4990 ;
      RECT 1.3430 0.4990 1.4330 0.5000 ;
      RECT 1.0390 0.5000 1.4330 0.5500 ;
      RECT 1.3830 0.5500 1.4330 0.6020 ;
      RECT 1.3430 0.9150 1.4330 0.9200 ;
      RECT 1.3430 0.9200 1.3930 1.1450 ;
      RECT 1.3830 0.6520 1.4330 0.8650 ;
      RECT 1.0390 0.8650 1.4330 0.9150 ;
      RECT 1.8330 0.1500 1.8830 0.3070 ;
      RECT 1.3430 0.3070 1.8830 0.3570 ;
      RECT 1.3830 0.6020 1.7890 0.6520 ;
      RECT 1.7470 1.5270 3.0050 1.5770 ;
      RECT 1.7470 1.2450 1.7970 1.5270 ;
      RECT 0.8870 1.1950 1.7970 1.2450 ;
      RECT 0.5830 0.8750 0.6330 1.5070 ;
      RECT 0.5830 0.1640 0.6330 0.4330 ;
      RECT 0.8870 1.2450 0.9370 1.5070 ;
      RECT 0.8870 0.8750 0.9370 1.1950 ;
      RECT 0.5830 0.8250 0.9770 0.8750 ;
      RECT 0.9270 0.4830 0.9770 0.8250 ;
      RECT 0.5830 0.4330 0.9770 0.4830 ;
      RECT 0.8870 0.1660 0.9370 0.4330 ;
      RECT 0.4860 0.6020 0.8770 0.6520 ;
      RECT 0.4310 0.7360 0.5360 0.7520 ;
      RECT 0.4310 0.7520 0.5350 0.7860 ;
      RECT 0.4310 0.1760 0.4810 0.5020 ;
      RECT 0.4310 0.7860 0.4810 1.2110 ;
      RECT 0.4860 0.6520 0.5360 0.7360 ;
      RECT 0.4860 0.5520 0.5360 0.6020 ;
      RECT 0.4310 0.5020 0.5360 0.5520 ;
      RECT 2.9220 0.6600 4.0840 0.7100 ;
      RECT 5.2430 0.5460 10.1640 0.5890 ;
      RECT 2.1030 0.5390 10.1640 0.5460 ;
      RECT 2.1030 0.3360 2.1530 0.4960 ;
      RECT 2.4070 0.3360 2.4570 0.4960 ;
      RECT 2.7110 0.3360 2.7610 0.4960 ;
      RECT 3.3190 0.3420 3.3690 0.4960 ;
      RECT 3.6230 0.3420 3.6730 0.4960 ;
      RECT 3.9270 0.3420 3.9770 0.4960 ;
      RECT 4.2310 0.3630 4.2810 0.4960 ;
      RECT 4.2310 0.8030 4.2810 1.1020 ;
      RECT 4.5350 0.3630 4.5850 0.4960 ;
      RECT 4.5350 0.8030 4.5850 1.1020 ;
      RECT 4.8390 0.3630 4.8890 0.4960 ;
      RECT 4.8390 0.8030 4.8890 1.1020 ;
      RECT 5.1430 0.5460 5.1930 0.7530 ;
      RECT 5.1430 0.3630 5.1930 0.4960 ;
      RECT 4.2310 0.7530 5.1930 0.8030 ;
      RECT 5.1430 0.8030 5.1930 0.9340 ;
      RECT 2.1030 0.4960 5.2930 0.5390 ;
  END
END TNBUFFX32_LVT

MACRO TNBUFFX4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.432 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3240 1.3730 0.7360 1.4230 ;
        RECT 0.5530 1.4230 0.6630 1.5750 ;
    END
    ANTENNAGATEAREA 0.0339 ;
  END EN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.4320 1.7020 ;
        RECT 1.9510 1.2720 2.0010 1.6420 ;
        RECT 1.6470 1.2750 1.6970 1.6420 ;
        RECT 0.2240 1.2560 0.2740 1.6420 ;
        RECT 0.8870 1.3210 0.9370 1.6420 ;
        RECT 0.2240 1.2060 0.3290 1.2560 ;
        RECT 0.7350 1.2710 0.9370 1.3210 ;
        RECT 0.2790 0.7310 0.3290 1.2060 ;
        RECT 0.7350 1.0900 0.7850 1.2710 ;
        RECT 0.8870 1.0900 0.9370 1.2710 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.4320 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.5420 ;
        RECT 1.9510 0.0300 2.0010 0.3680 ;
        RECT 1.6470 0.0300 1.6970 0.1910 ;
        RECT 1.0390 0.1910 1.6970 0.2410 ;
        RECT 1.0390 0.2410 1.0890 0.4530 ;
        RECT 1.1920 0.2410 1.2420 0.4530 ;
        RECT 1.6470 0.2410 1.6970 0.3680 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4950 0.4380 2.2150 0.4880 ;
        RECT 2.1650 0.4880 2.3350 0.6630 ;
        RECT 2.1030 0.1550 2.1530 0.4380 ;
        RECT 1.7990 0.1420 1.8490 0.4380 ;
        RECT 1.4950 0.2910 1.5450 0.4380 ;
        RECT 2.1650 0.6630 2.2150 1.0840 ;
        RECT 1.4950 1.0840 2.2150 1.1340 ;
        RECT 2.1030 1.1340 2.1530 1.4720 ;
        RECT 1.7990 1.1340 1.8490 1.4720 ;
        RECT 1.7990 0.9000 1.8490 1.0840 ;
        RECT 1.4950 1.1340 1.5450 1.4720 ;
    END
    ANTENNADIFFAREA 0.3552 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 0.6460 1.0440 0.6960 ;
        RECT 0.8570 0.6960 0.9670 0.8150 ;
    END
    ANTENNAGATEAREA 0.0366 ;
  END A
  OBS
    LAYER NWELL ;
      RECT -0.1120 0.6790 2.5440 1.7730 ;
    LAYER M1 ;
      RECT 0.8870 0.5390 2.1050 0.5890 ;
      RECT 0.8870 0.5890 0.9370 0.5900 ;
      RECT 0.8870 0.4890 0.9370 0.5390 ;
      RECT 0.7350 0.4390 0.9370 0.4890 ;
      RECT 0.8870 0.2550 0.9370 0.4390 ;
      RECT 1.3430 0.5890 1.3930 0.9340 ;
      RECT 1.3430 0.2910 1.3930 0.5390 ;
      RECT 0.7350 0.2550 0.7850 0.4390 ;
      RECT 1.5400 0.7450 2.1080 0.7950 ;
      RECT 1.0390 1.0340 1.0890 1.4780 ;
      RECT 1.0390 0.8050 1.0890 0.9840 ;
      RECT 1.1920 1.0340 1.2420 1.2020 ;
      RECT 1.1920 0.7130 1.2420 0.9840 ;
      RECT 0.5830 0.1910 0.6330 0.9840 ;
      RECT 0.5830 1.0340 0.6330 1.3230 ;
      RECT 1.5710 0.7950 1.6210 0.9840 ;
      RECT 0.5830 0.9840 1.6210 1.0340 ;
      RECT 0.4310 0.0910 1.3480 0.1410 ;
      RECT 0.4310 0.1410 0.4810 1.2110 ;
    LAYER PO ;
      RECT 1.7330 0.7170 1.7630 1.6060 ;
      RECT 1.8850 0.7170 1.9150 1.6060 ;
      RECT 2.0370 0.7170 2.0670 1.6060 ;
      RECT 1.5810 0.7170 1.6110 1.6060 ;
      RECT 1.5810 0.0660 1.6110 0.6170 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 2.0370 0.0660 2.0670 0.6170 ;
      RECT 1.8850 0.0660 1.9150 0.6170 ;
      RECT 1.7330 0.0660 1.7630 0.6170 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
  END
END TNBUFFX4_LVT

MACRO TNBUFFX8_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.496 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3240 1.3730 0.8880 1.4230 ;
        RECT 0.7050 1.4230 0.8150 1.5750 ;
    END
    ANTENNAGATEAREA 0.0522 ;
  END EN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.4960 1.7020 ;
        RECT 3.0150 1.2720 3.0650 1.6420 ;
        RECT 2.7110 1.2720 2.7610 1.6420 ;
        RECT 2.4070 1.2720 2.4570 1.6420 ;
        RECT 2.1030 1.2750 2.1530 1.6420 ;
        RECT 0.2240 1.2560 0.2740 1.6420 ;
        RECT 1.1910 1.3210 1.2410 1.6420 ;
        RECT 0.2240 1.2060 0.3290 1.2560 ;
        RECT 0.5830 1.2710 1.2410 1.3210 ;
        RECT 0.2790 0.7310 0.3290 1.2060 ;
        RECT 0.5830 0.8140 0.6330 1.2710 ;
        RECT 0.8870 1.0840 0.9370 1.2710 ;
        RECT 1.1910 1.0840 1.2410 1.2710 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.4960 0.0300 ;
        RECT 3.0150 0.0300 3.0650 0.3680 ;
        RECT 2.7110 0.0300 2.7610 0.3680 ;
        RECT 0.2790 0.0300 0.3290 0.5740 ;
        RECT 2.4070 0.0300 2.4570 0.3680 ;
        RECT 2.1030 0.0300 2.1530 0.1910 ;
        RECT 1.0390 0.1910 2.1530 0.2410 ;
        RECT 1.3430 0.2410 1.3930 0.4360 ;
        RECT 1.6480 0.2410 1.6980 0.4880 ;
        RECT 1.0390 0.2410 1.0890 0.3950 ;
        RECT 2.1030 0.2410 2.1530 0.3680 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2290 0.4890 3.2790 0.6370 ;
        RECT 3.2290 0.6370 3.4260 0.8150 ;
        RECT 3.1670 0.4880 3.2790 0.4890 ;
        RECT 3.2290 0.8150 3.2790 1.0840 ;
        RECT 1.9510 0.4390 3.2790 0.4880 ;
        RECT 1.9510 1.0840 3.2790 1.1340 ;
        RECT 1.9510 0.4380 3.2410 0.4390 ;
        RECT 3.1670 1.1340 3.2170 1.4720 ;
        RECT 2.8630 1.1340 2.9130 1.4720 ;
        RECT 2.8630 0.9000 2.9130 1.0840 ;
        RECT 2.5590 1.1340 2.6090 1.4720 ;
        RECT 2.5590 0.9000 2.6090 1.0840 ;
        RECT 2.2550 1.1340 2.3050 1.4720 ;
        RECT 2.2550 0.9000 2.3050 1.0840 ;
        RECT 1.9510 1.1340 2.0010 1.4720 ;
        RECT 3.1670 0.1550 3.2170 0.4380 ;
        RECT 2.8630 0.1420 2.9130 0.4380 ;
        RECT 2.5590 0.1420 2.6090 0.4380 ;
        RECT 2.2550 0.1420 2.3050 0.4380 ;
        RECT 1.9510 0.2910 2.0010 0.4380 ;
    END
    ANTENNADIFFAREA 0.6212 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0090 0.6600 1.3480 0.7100 ;
        RECT 1.0090 0.7100 1.1190 0.8150 ;
    END
    ANTENNAGATEAREA 0.0732 ;
  END A
  OBS
    LAYER NWELL ;
      RECT -0.1120 0.6790 3.6110 1.7730 ;
    LAYER M1 ;
      RECT 0.8870 0.5390 3.1720 0.5770 ;
      RECT 0.8870 0.5770 3.1690 0.5890 ;
      RECT 1.1910 0.3280 1.2410 0.5390 ;
      RECT 1.4950 0.3480 1.5450 0.5390 ;
      RECT 1.7990 0.3480 1.8490 0.5390 ;
      RECT 1.7990 0.5890 1.8490 0.8840 ;
      RECT 1.4640 0.8840 1.8490 0.9340 ;
      RECT 0.8870 0.2410 0.9370 0.5390 ;
      RECT 0.5830 0.1910 0.9370 0.2410 ;
      RECT 0.5830 0.2410 0.6330 0.4870 ;
      RECT 1.9960 0.7450 3.1690 0.7950 ;
      RECT 1.0390 1.0340 1.0890 1.2020 ;
      RECT 1.0390 0.9060 1.0890 0.9840 ;
      RECT 1.3430 1.0340 1.3930 1.4780 ;
      RECT 1.3430 0.8140 1.3930 0.9840 ;
      RECT 1.6480 1.0340 1.6980 1.2940 ;
      RECT 0.7350 1.0340 0.7850 1.1190 ;
      RECT 0.7350 0.3750 0.7850 0.9840 ;
      RECT 2.0270 0.7950 2.0770 0.9840 ;
      RECT 0.7350 0.9840 2.0770 1.0340 ;
      RECT 0.4310 0.0910 1.8040 0.1410 ;
      RECT 0.4310 0.1410 0.4810 1.2110 ;
    LAYER PO ;
      RECT 2.4930 0.0660 2.5230 0.6170 ;
      RECT 2.3410 0.0660 2.3710 0.6170 ;
      RECT 2.1890 0.0660 2.2190 0.6170 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 2.7970 0.0660 2.8270 0.6170 ;
      RECT 2.7970 0.7170 2.8270 1.6060 ;
      RECT 3.1010 0.0660 3.1310 0.6170 ;
      RECT 3.1010 0.7170 3.1310 1.6060 ;
      RECT 2.9490 0.0660 2.9790 0.6170 ;
      RECT 2.9490 0.7170 2.9790 1.6060 ;
      RECT 2.6450 0.0660 2.6750 0.6170 ;
      RECT 2.6450 0.7170 2.6750 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 2.1890 0.7170 2.2190 1.6060 ;
      RECT 2.3410 0.7170 2.3710 1.6060 ;
      RECT 2.4930 0.7170 2.5230 1.6060 ;
      RECT 2.0370 0.7170 2.0670 1.6060 ;
      RECT 2.0370 0.0660 2.0670 0.6170 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
  END
END TNBUFFX8_LVT

MACRO XNOR2X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.584 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.5840 1.7020 ;
        RECT 1.0390 1.2180 1.0890 1.6420 ;
        RECT 0.2790 1.1290 0.3290 1.6420 ;
        RECT 2.1030 0.8140 2.1530 1.6420 ;
        RECT 1.6470 1.2180 1.6970 1.6420 ;
        RECT 0.5830 1.2180 0.6330 1.6420 ;
    END
  END VDD

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6580 0.7050 0.8150 0.8030 ;
        RECT 0.6580 0.8030 1.6550 0.8530 ;
    END
    ANTENNAGATEAREA 0.0378 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9620 0.6720 1.9410 0.7220 ;
        RECT 0.9620 0.5530 1.1190 0.6720 ;
    END
    ANTENNAGATEAREA 0.0405 ;
  END A1

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.5840 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.3710 ;
        RECT 2.1030 0.0300 2.1530 0.5260 ;
        RECT 1.7350 0.0300 1.7850 0.2700 ;
        RECT 0.2790 0.3710 0.6120 0.4210 ;
        RECT 1.6160 0.2700 1.7850 0.3200 ;
        RECT 0.5620 0.3200 0.6120 0.3710 ;
        RECT 0.5620 0.2700 1.1200 0.3200 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2550 0.9170 2.4870 0.9670 ;
        RECT 2.3100 0.8570 2.4870 0.9170 ;
        RECT 2.2550 0.9670 2.3050 1.5460 ;
        RECT 2.3100 0.5540 2.3600 0.8570 ;
        RECT 2.2550 0.5040 2.3600 0.5540 ;
        RECT 2.2550 0.1480 2.3050 0.5040 ;
    END
    ANTENNADIFFAREA 0.1234 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 2.6990 1.7810 ;
    LAYER M1 ;
      RECT 0.3550 1.0180 0.8160 1.0680 ;
      RECT 0.7350 0.3700 0.7850 0.4710 ;
      RECT 0.3550 0.6540 0.4050 1.0180 ;
      RECT 0.3240 0.6040 0.4050 0.6540 ;
      RECT 0.3550 0.5210 0.4050 0.6040 ;
      RECT 0.3550 0.4710 0.7850 0.5210 ;
      RECT 0.8460 0.4080 1.2240 0.4580 ;
      RECT 1.1740 0.4580 1.2240 0.5720 ;
      RECT 0.4800 0.9180 0.9370 0.9680 ;
      RECT 0.8870 0.9680 0.9370 1.0680 ;
      RECT 1.1740 0.5720 1.3500 0.6220 ;
      RECT 0.8460 0.4580 0.8960 0.5710 ;
      RECT 0.4800 0.5710 0.8960 0.6210 ;
      RECT 0.4800 0.6210 0.5300 0.9180 ;
      RECT 1.9910 0.6040 2.2600 0.6540 ;
      RECT 1.3600 0.3750 1.4100 0.4710 ;
      RECT 1.3270 0.3250 1.4100 0.3750 ;
      RECT 1.9910 0.5210 2.0410 0.6040 ;
      RECT 1.9510 0.8090 2.0410 0.8590 ;
      RECT 1.3600 0.4710 2.0410 0.5210 ;
      RECT 1.9510 0.8590 2.0010 1.0080 ;
      RECT 1.9510 0.2400 2.0010 0.4710 ;
      RECT 1.3120 1.0080 2.0010 1.0580 ;
      RECT 1.9510 1.0580 2.0010 1.3050 ;
      RECT 1.9910 0.6540 2.0410 0.8090 ;
      RECT 0.4620 0.1530 1.2410 0.2030 ;
      RECT 1.1910 0.2030 1.2410 0.3260 ;
      RECT 0.4620 0.2030 0.5120 0.2710 ;
      RECT 0.4000 0.2710 0.5120 0.3210 ;
      RECT 1.4640 0.3710 1.8800 0.4210 ;
      RECT 1.1600 1.2390 1.5760 1.2890 ;
      RECT 1.7990 1.1680 1.8490 1.3200 ;
      RECT 0.4310 1.1180 1.8490 1.1680 ;
      RECT 0.4310 1.1680 0.4810 1.3200 ;
    LAYER PO ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 1.2770 0.0680 1.3070 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
  END
END XNOR2X1_LVT

MACRO XNOR2X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.736 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6580 0.8030 1.6210 0.8530 ;
        RECT 0.6580 0.6440 0.8150 0.8030 ;
        RECT 1.5710 0.6270 1.6210 0.8030 ;
    END
    ANTENNAGATEAREA 0.066 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4190 0.4690 1.9250 0.5190 ;
        RECT 1.8750 0.5190 1.9250 0.6530 ;
        RECT 1.4190 0.5190 1.4690 0.6720 ;
        RECT 0.9620 0.6720 1.4690 0.7220 ;
        RECT 0.9620 0.5530 1.1190 0.6720 ;
    END
    ANTENNAGATEAREA 0.0708 ;
  END A1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.7360 1.7020 ;
        RECT 2.4070 1.0750 2.4570 1.6420 ;
        RECT 2.1030 0.8140 2.1530 1.6420 ;
        RECT 0.2790 1.1930 0.3290 1.6420 ;
        RECT 1.0390 1.2850 1.0890 1.6420 ;
        RECT 1.6470 1.2850 1.6970 1.6420 ;
        RECT 0.5830 1.2850 0.6330 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.7360 0.0300 ;
        RECT 2.1030 0.0300 2.1530 0.5200 ;
        RECT 2.4070 0.0300 2.4570 0.4160 ;
        RECT 0.2790 0.0300 0.3290 0.1630 ;
        RECT 1.6940 0.0300 1.7440 0.1620 ;
        RECT 0.2790 0.1630 1.1200 0.2130 ;
        RECT 1.6180 0.1620 1.7440 0.2120 ;
        RECT 0.2790 0.2130 0.3290 0.2380 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2550 0.9340 2.5220 0.9840 ;
        RECT 2.2550 0.9840 2.3050 1.5460 ;
        RECT 2.3770 0.8570 2.5220 0.9340 ;
        RECT 2.4720 0.5540 2.5220 0.8570 ;
        RECT 2.2550 0.5040 2.5220 0.5540 ;
        RECT 2.2550 0.1480 2.3050 0.5040 ;
    END
    ANTENNADIFFAREA 0.1464 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 2.8510 1.7810 ;
    LAYER M1 ;
      RECT 0.3240 1.0180 0.8160 1.0680 ;
      RECT 0.3240 0.3630 0.8010 0.4130 ;
      RECT 0.3240 0.6540 0.3740 1.0180 ;
      RECT 0.3240 0.6040 0.4210 0.6540 ;
      RECT 0.3240 0.4130 0.3740 0.6040 ;
      RECT 0.8710 0.4080 1.2240 0.4580 ;
      RECT 1.1740 0.4580 1.2240 0.5720 ;
      RECT 0.8710 0.4580 0.9210 0.4630 ;
      RECT 0.4800 0.9180 0.9530 0.9680 ;
      RECT 1.1740 0.5720 1.3500 0.6220 ;
      RECT 0.4800 0.4630 0.9210 0.5030 ;
      RECT 0.4800 0.5030 0.9120 0.5130 ;
      RECT 0.4800 0.5130 0.5300 0.9180 ;
      RECT 1.9890 0.6040 2.4140 0.6540 ;
      RECT 1.9890 0.6540 2.0390 0.8090 ;
      RECT 1.9890 0.4120 2.0390 0.6040 ;
      RECT 1.9510 0.8090 2.0390 0.8590 ;
      RECT 1.3070 0.3620 2.0390 0.4120 ;
      RECT 1.9510 0.8590 2.0010 1.0080 ;
      RECT 1.9510 0.2400 2.0010 0.3620 ;
      RECT 1.3120 1.0080 2.0010 1.0580 ;
      RECT 1.9510 1.0580 2.0010 1.5550 ;
      RECT 1.4640 0.2620 1.8800 0.3120 ;
      RECT 1.1600 1.2390 1.5760 1.2890 ;
      RECT 0.4310 1.1180 1.8490 1.1680 ;
      RECT 1.7990 1.1680 1.8490 1.3200 ;
      RECT 0.4310 1.1680 0.4810 1.5510 ;
      RECT 0.4010 0.2630 1.2570 0.3130 ;
    LAYER PO ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 1.2770 0.0680 1.3070 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
  END
END XNOR2X2_LVT

MACRO XNOR3X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.648 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4670 0.1160 2.6200 0.1660 ;
        RECT 2.5700 0.1660 2.6200 0.3500 ;
        RECT 2.5700 0.3500 2.7560 0.4000 ;
        RECT 2.7060 0.4000 2.7560 0.6190 ;
        RECT 2.7060 0.6190 2.9900 0.6690 ;
        RECT 2.8330 0.5530 2.9900 0.6190 ;
    END
    ANTENNAGATEAREA 0.0465 ;
  END A3

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.3190 0.4620 3.5510 0.5120 ;
        RECT 3.3990 0.5120 3.4490 0.8020 ;
        RECT 3.3190 0.1280 3.3690 0.4620 ;
        RECT 3.4330 0.4010 3.5510 0.4620 ;
        RECT 3.3190 0.8020 3.4490 0.8520 ;
        RECT 3.3190 0.8520 3.3690 1.5460 ;
    END
    ANTENNADIFFAREA 0.1142 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.6480 1.7020 ;
        RECT 1.6470 1.3050 1.6970 1.6420 ;
        RECT 0.2790 0.9440 0.3290 1.6420 ;
        RECT 2.1030 1.2150 2.1530 1.6420 ;
        RECT 3.1670 1.2990 3.2170 1.6420 ;
        RECT 0.5830 1.3710 0.6330 1.6420 ;
        RECT 2.8470 1.2490 3.2170 1.2990 ;
        RECT 0.5830 1.3210 1.1050 1.3710 ;
        RECT 0.5830 1.3040 0.6330 1.3210 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.6480 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.3910 ;
        RECT 2.1030 0.0300 2.1530 0.3430 ;
        RECT 1.7350 0.0300 1.7850 0.2340 ;
        RECT 3.1670 0.0300 3.2170 0.2740 ;
        RECT 0.2790 0.3910 0.5810 0.4410 ;
        RECT 1.6310 0.2340 1.7850 0.2840 ;
        RECT 2.8470 0.2740 3.2170 0.3240 ;
        RECT 0.5310 0.3200 0.5810 0.3910 ;
        RECT 0.5310 0.2700 1.1050 0.3200 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9620 1.4650 1.1190 1.5750 ;
    END
    ANTENNAGATEAREA 0.057 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6600 0.7050 0.8150 0.8260 ;
        RECT 0.6600 0.8260 1.6210 0.8760 ;
        RECT 1.5710 0.7030 1.6210 0.8260 ;
    END
    ANTENNAGATEAREA 0.0555 ;
  END A2
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 3.7630 1.7810 ;
    LAYER M1 ;
      RECT 1.4180 0.5340 1.9250 0.5840 ;
      RECT 1.8750 0.5840 1.9250 0.7540 ;
      RECT 1.4180 0.5840 1.4680 0.7030 ;
      RECT 0.9470 0.7030 1.4680 0.7530 ;
      RECT 2.6870 1.4850 2.8530 1.5350 ;
      RECT 1.9510 1.1650 2.0010 1.3770 ;
      RECT 1.3270 1.1040 2.0010 1.1150 ;
      RECT 1.9510 0.8590 2.0010 1.1040 ;
      RECT 1.9510 0.2440 2.0010 0.4340 ;
      RECT 2.6870 1.2990 2.7370 1.4850 ;
      RECT 2.3580 1.2490 2.7370 1.2990 ;
      RECT 2.3580 1.1650 2.4080 1.2490 ;
      RECT 1.3270 1.1150 2.4080 1.1540 ;
      RECT 1.9510 0.8090 2.2450 0.8590 ;
      RECT 2.0060 0.4840 2.0560 0.8090 ;
      RECT 1.3590 0.4340 2.0560 0.4840 ;
      RECT 1.9510 1.1540 2.4080 1.1650 ;
      RECT 1.3590 0.3750 1.4090 0.4340 ;
      RECT 1.3260 0.3250 1.4090 0.3750 ;
      RECT 0.4340 1.0990 0.8010 1.1490 ;
      RECT 0.7350 0.3770 0.7850 0.4910 ;
      RECT 0.4340 0.4910 0.7850 0.5410 ;
      RECT 0.4340 0.6540 0.4840 1.0990 ;
      RECT 0.3390 0.6040 0.4840 0.6540 ;
      RECT 0.4340 0.5410 0.4840 0.6040 ;
      RECT 0.5490 0.9990 0.9530 1.0490 ;
      RECT 0.5490 0.5910 0.8880 0.6410 ;
      RECT 0.8380 0.4580 0.8880 0.5910 ;
      RECT 0.8380 0.4080 1.2360 0.4580 ;
      RECT 1.1860 0.4580 1.2360 0.5930 ;
      RECT 1.1860 0.5930 1.3500 0.6430 ;
      RECT 0.5490 0.6410 0.5990 0.9990 ;
      RECT 0.4310 1.2040 1.8650 1.2540 ;
      RECT 0.4310 1.2540 0.4810 1.3200 ;
      RECT 2.7110 0.1110 2.8530 0.1610 ;
      RECT 2.7110 0.1610 2.7610 0.3000 ;
      RECT 3.1570 0.6040 3.3090 0.6540 ;
      RECT 3.1570 0.6540 3.2070 1.1490 ;
      RECT 2.5430 1.1490 3.2070 1.1990 ;
      RECT 2.8340 0.8720 2.8840 1.1490 ;
      RECT 2.3950 0.8220 2.8840 0.8720 ;
      RECT 2.3950 0.5000 2.4450 0.8220 ;
      RECT 2.3950 0.4500 2.6250 0.5000 ;
      RECT 0.4310 0.1530 1.2410 0.2030 ;
      RECT 1.1910 0.2030 1.2410 0.3000 ;
      RECT 0.4310 0.2030 0.4810 0.3410 ;
      RECT 2.9990 0.9890 3.0900 1.0390 ;
      RECT 3.0400 0.7690 3.0900 0.9890 ;
      RECT 2.9990 0.3740 3.0900 0.4240 ;
      RECT 2.6040 0.7190 3.0900 0.7690 ;
      RECT 3.0400 0.4240 3.0900 0.7190 ;
      RECT 2.2380 0.9840 2.7770 1.0340 ;
      RECT 2.2950 0.2970 2.3450 0.9840 ;
      RECT 2.2390 0.2470 2.4730 0.2970 ;
      RECT 1.4790 0.3340 1.8650 0.3840 ;
      RECT 1.1750 1.3210 1.5610 1.3710 ;
    LAYER PO ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 1.2770 0.0680 1.3070 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
  END
END XNOR3X1_LVT

MACRO XNOR3X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9620 1.4650 1.1190 1.5750 ;
    END
    ANTENNAGATEAREA 0.0531 ;
  END A1

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.7060 0.4100 2.7560 0.6190 ;
        RECT 2.7060 0.6190 2.9910 0.6690 ;
        RECT 2.5700 0.3600 2.7560 0.4100 ;
        RECT 2.8330 0.5530 2.9900 0.6190 ;
        RECT 2.5700 0.1640 2.6200 0.3600 ;
        RECT 2.4670 0.1140 2.6200 0.1640 ;
    END
    ANTENNAGATEAREA 0.0504 ;
  END A3

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.8000 1.7020 ;
        RECT 3.4710 0.9210 3.5210 1.6420 ;
        RECT 1.6470 1.2430 1.6970 1.6420 ;
        RECT 0.2790 0.9440 0.3290 1.6420 ;
        RECT 2.1030 1.2150 2.1530 1.6420 ;
        RECT 3.1670 1.2990 3.2170 1.6420 ;
        RECT 0.5830 1.3090 0.6330 1.6420 ;
        RECT 2.8470 1.2490 3.2170 1.2990 ;
        RECT 0.5830 1.2590 1.1050 1.3090 ;
        RECT 0.5830 1.2420 0.6330 1.2590 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.8000 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.3910 ;
        RECT 3.4710 0.0300 3.5210 0.3190 ;
        RECT 2.1030 0.0300 2.1530 0.3430 ;
        RECT 1.6470 0.0300 1.6970 0.2730 ;
        RECT 3.1670 0.0300 3.2170 0.2580 ;
        RECT 0.2790 0.3910 0.5810 0.4410 ;
        RECT 2.8470 0.2580 3.2170 0.3080 ;
        RECT 0.5310 0.3200 0.5810 0.3910 ;
        RECT 3.1670 0.3080 3.2170 0.3240 ;
        RECT 0.5310 0.2700 1.1200 0.3200 ;
    END
  END VSS

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6600 0.7050 0.8150 0.8260 ;
        RECT 0.6600 0.8260 1.6210 0.8760 ;
        RECT 1.5710 0.7030 1.6210 0.8260 ;
    END
    ANTENNAGATEAREA 0.0531 ;
  END A2

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4410 0.4010 3.5510 0.5040 ;
        RECT 3.3190 0.5040 3.5610 0.5540 ;
        RECT 3.3190 0.1480 3.3690 0.5040 ;
        RECT 3.5110 0.5540 3.5610 0.7820 ;
        RECT 3.3190 0.7820 3.5610 0.8320 ;
        RECT 3.3190 0.8320 3.3690 1.5460 ;
    END
    ANTENNADIFFAREA 0.1464 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 3.9150 1.7810 ;
    LAYER M1 ;
      RECT 1.4180 0.5340 1.9250 0.5840 ;
      RECT 1.8750 0.5840 1.9250 0.7540 ;
      RECT 1.4180 0.5840 1.4680 0.7030 ;
      RECT 0.9470 0.7030 1.4680 0.7530 ;
      RECT 2.5420 1.0890 3.2690 1.1390 ;
      RECT 3.2190 0.6540 3.2690 1.0890 ;
      RECT 3.2190 0.6040 3.4610 0.6540 ;
      RECT 2.8790 0.8720 2.9290 1.0890 ;
      RECT 2.4290 0.8220 2.9290 0.8720 ;
      RECT 2.4290 0.5420 2.4790 0.8220 ;
      RECT 2.4290 0.4920 2.6250 0.5420 ;
      RECT 2.6870 1.4620 2.8530 1.5120 ;
      RECT 1.9510 1.1650 2.0010 1.3150 ;
      RECT 1.9510 1.0870 2.0010 1.1150 ;
      RECT 1.3120 1.0370 2.0010 1.0870 ;
      RECT 1.9510 0.8590 2.0010 1.0370 ;
      RECT 1.9510 0.2030 2.0010 0.4340 ;
      RECT 2.6870 1.2720 2.7370 1.4620 ;
      RECT 2.3910 1.2220 2.7370 1.2720 ;
      RECT 1.9510 0.8090 2.0560 0.8590 ;
      RECT 2.0060 0.6540 2.0560 0.8090 ;
      RECT 2.0060 0.6040 2.2450 0.6540 ;
      RECT 2.0060 0.4840 2.0560 0.6040 ;
      RECT 1.3610 0.4340 2.0560 0.4840 ;
      RECT 2.3910 1.1650 2.4410 1.2220 ;
      RECT 1.9510 1.1150 2.4410 1.1650 ;
      RECT 1.3610 0.3750 1.4110 0.4340 ;
      RECT 1.3270 0.3250 1.4110 0.3750 ;
      RECT 0.3900 1.0370 0.8160 1.0870 ;
      RECT 0.7350 0.3770 0.7850 0.4910 ;
      RECT 0.3900 0.4910 0.7850 0.5410 ;
      RECT 0.3900 0.6540 0.4400 1.0370 ;
      RECT 0.3240 0.6040 0.4400 0.6540 ;
      RECT 0.3900 0.5410 0.4400 0.6040 ;
      RECT 0.5280 0.9370 0.9530 0.9870 ;
      RECT 0.5280 0.5910 0.9020 0.6410 ;
      RECT 0.8520 0.4580 0.9020 0.5910 ;
      RECT 0.8520 0.4080 1.2440 0.4580 ;
      RECT 1.1940 0.4580 1.2440 0.5930 ;
      RECT 1.1940 0.5930 1.3500 0.6430 ;
      RECT 0.5280 0.6410 0.5780 0.9370 ;
      RECT 1.1600 1.2590 1.5760 1.3090 ;
      RECT 0.4310 1.1370 1.8490 1.1870 ;
      RECT 1.7990 1.1870 1.8490 1.2530 ;
      RECT 0.4310 1.1870 0.4810 1.2530 ;
      RECT 2.2190 0.9290 2.7770 0.9790 ;
      RECT 2.2950 0.2970 2.3450 0.9290 ;
      RECT 2.2390 0.2470 2.4880 0.2970 ;
      RECT 0.4310 0.1530 1.2410 0.2030 ;
      RECT 1.1910 0.2030 1.2410 0.3080 ;
      RECT 0.4310 0.2030 0.4810 0.3410 ;
      RECT 2.9980 0.9210 3.1270 0.9710 ;
      RECT 3.0770 0.7690 3.1270 0.9210 ;
      RECT 3.0770 0.4680 3.1270 0.7190 ;
      RECT 2.9840 0.4180 3.1270 0.4680 ;
      RECT 2.6190 0.7190 3.1270 0.7690 ;
      RECT 1.4790 0.3340 1.8700 0.3840 ;
      RECT 2.7110 0.1110 2.8530 0.1610 ;
      RECT 2.7110 0.1610 2.7610 0.2730 ;
    LAYER PO ;
      RECT 3.7090 0.0680 3.7390 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 1.2770 0.0680 1.3070 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
  END
END XNOR3X2_LVT

MACRO XOR2X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.584 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2550 0.7650 2.4870 0.8150 ;
        RECT 2.3100 0.7050 2.4870 0.7650 ;
        RECT 2.2550 0.8150 2.3050 1.5460 ;
        RECT 2.3100 0.5540 2.3600 0.7050 ;
        RECT 2.2550 0.5040 2.3600 0.5540 ;
        RECT 2.2550 0.1480 2.3050 0.5040 ;
    END
    ANTENNADIFFAREA 0.1193 ;
  END Y

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4000 0.7050 1.6520 0.7550 ;
        RECT 1.4000 0.7550 1.4500 0.7810 ;
        RECT 0.5530 0.7810 1.4500 0.8150 ;
        RECT 0.5530 0.7050 0.7110 0.7810 ;
        RECT 0.5550 0.8150 1.4500 0.8310 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 0.5530 1.0510 0.6630 ;
        RECT 1.0010 0.6630 1.0510 0.6710 ;
        RECT 1.0010 0.6710 1.3480 0.7210 ;
    END
    ANTENNAGATEAREA 0.0336 ;
  END A1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.5840 1.7020 ;
        RECT 0.2790 0.9440 0.3290 1.6420 ;
        RECT 1.6470 1.2080 1.6970 1.6420 ;
        RECT 0.5830 1.2080 0.6330 1.6420 ;
        RECT 1.0390 1.2080 1.0890 1.6420 ;
        RECT 2.1030 0.8140 2.1530 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.5840 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.4020 ;
        RECT 2.1030 0.0300 2.1530 0.0980 ;
        RECT 0.2790 0.4020 0.5960 0.4520 ;
        RECT 1.7350 0.0980 2.1530 0.1480 ;
        RECT 0.5460 0.3500 0.5960 0.4020 ;
        RECT 1.7350 0.1480 1.7850 0.2700 ;
        RECT 2.1030 0.1480 2.1530 0.4280 ;
        RECT 0.5460 0.3000 1.1200 0.3500 ;
        RECT 1.6160 0.2700 1.7850 0.3200 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 2.6990 1.7810 ;
    LAYER M1 ;
      RECT 0.4030 0.5190 0.7850 0.5690 ;
      RECT 0.7350 0.4020 0.7850 0.5190 ;
      RECT 0.4030 1.0080 0.8010 1.0580 ;
      RECT 0.4030 0.5690 0.4530 0.6040 ;
      RECT 0.3240 0.6040 0.4530 0.6540 ;
      RECT 0.4030 0.6540 0.4530 1.0080 ;
      RECT 1.7990 1.1580 1.8490 1.3200 ;
      RECT 0.4310 1.1080 1.8490 1.1580 ;
      RECT 0.4310 1.1580 0.4810 1.3200 ;
      RECT 1.1130 0.8900 1.7520 0.9400 ;
      RECT 1.7020 0.6210 1.7520 0.8900 ;
      RECT 1.1700 0.4580 1.2200 0.5710 ;
      RECT 0.8710 0.4080 1.2200 0.4580 ;
      RECT 1.1130 0.9400 1.1630 1.0080 ;
      RECT 0.8710 1.0080 1.1630 1.0580 ;
      RECT 1.1700 0.5710 1.9560 0.6210 ;
      RECT 2.0060 0.6040 2.2600 0.6540 ;
      RECT 2.0060 0.6540 2.0560 0.7040 ;
      RECT 2.0060 0.5210 2.0560 0.6040 ;
      RECT 1.9510 0.7040 2.0560 0.7540 ;
      RECT 1.3430 0.4780 2.0560 0.5210 ;
      RECT 1.3430 0.4710 2.0530 0.4780 ;
      RECT 1.3430 0.2940 1.3930 0.4710 ;
      RECT 1.9510 0.7540 2.0010 1.0080 ;
      RECT 1.9510 0.2400 2.0010 0.4710 ;
      RECT 1.3120 1.0080 2.0010 1.0580 ;
      RECT 1.9510 1.0580 2.0010 1.3150 ;
      RECT 1.1600 1.2390 1.5760 1.2890 ;
      RECT 1.4640 0.3710 1.8800 0.4210 ;
      RECT 0.4310 0.1530 1.2410 0.2030 ;
      RECT 1.1910 0.2030 1.2410 0.3260 ;
      RECT 0.4310 0.2030 0.4810 0.3520 ;
    LAYER PO ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 1.2770 0.0680 1.3070 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
  END
END XOR2X1_LVT

MACRO XOR2X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.736 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2540 0.7820 2.4970 0.8320 ;
        RECT 2.2540 0.8320 2.3040 1.5460 ;
        RECT 2.3770 0.7050 2.4970 0.7820 ;
        RECT 2.4470 0.5500 2.4970 0.7050 ;
        RECT 2.2540 0.5000 2.4970 0.5500 ;
        RECT 2.2540 0.1480 2.3040 0.5000 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 0.5530 1.0510 0.6630 ;
        RECT 1.0010 0.6630 1.0510 0.6710 ;
        RECT 1.0010 0.6710 1.3480 0.7210 ;
    END
    ANTENNAGATEAREA 0.0594 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4000 0.7050 1.6520 0.7550 ;
        RECT 1.4000 0.7550 1.4500 0.7810 ;
        RECT 0.5530 0.7810 1.4500 0.8150 ;
        RECT 0.5530 0.7050 0.7110 0.7810 ;
        RECT 0.5550 0.8150 1.4500 0.8310 ;
    END
    ANTENNAGATEAREA 0.0606 ;
  END A2

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.7360 1.7020 ;
        RECT 2.1030 0.8140 2.1530 1.6420 ;
        RECT 2.4070 0.9740 2.4570 1.6420 ;
        RECT 0.2790 0.9440 0.3290 1.6420 ;
        RECT 1.0390 1.2080 1.0890 1.6420 ;
        RECT 1.6470 1.2080 1.6970 1.6420 ;
        RECT 0.5830 1.2080 0.6330 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.7360 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.4020 ;
        RECT 2.4070 0.0300 2.4570 0.4370 ;
        RECT 2.1030 0.0300 2.1530 0.0980 ;
        RECT 0.2790 0.4020 0.5960 0.4520 ;
        RECT 1.7350 0.0980 2.1530 0.1480 ;
        RECT 0.5460 0.3200 0.5960 0.4020 ;
        RECT 1.7350 0.1480 1.7850 0.2700 ;
        RECT 2.1030 0.1480 2.1530 0.4160 ;
        RECT 0.5460 0.2700 1.1200 0.3200 ;
        RECT 1.6160 0.2700 1.7850 0.3200 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 2.8510 1.7810 ;
    LAYER M1 ;
      RECT 0.4030 1.0080 0.8010 1.0580 ;
      RECT 0.4030 0.5190 0.7850 0.5690 ;
      RECT 0.7350 0.3770 0.7850 0.5190 ;
      RECT 0.4030 0.6540 0.4530 1.0080 ;
      RECT 0.3240 0.6040 0.4530 0.6540 ;
      RECT 0.4030 0.5690 0.4530 0.6040 ;
      RECT 2.0060 0.6040 2.3970 0.6540 ;
      RECT 1.3430 0.2940 1.3930 0.4710 ;
      RECT 1.9510 0.2400 2.0010 0.4710 ;
      RECT 1.9510 0.7540 2.0010 1.0080 ;
      RECT 1.3120 1.0080 2.0010 1.0580 ;
      RECT 1.9510 1.0580 2.0010 1.3150 ;
      RECT 2.0060 0.5210 2.0560 0.6040 ;
      RECT 2.0060 0.6540 2.0560 0.7040 ;
      RECT 1.3430 0.4710 2.0560 0.5210 ;
      RECT 1.9510 0.7040 2.0560 0.7540 ;
      RECT 1.1600 1.2390 1.5760 1.2890 ;
      RECT 1.1130 0.8900 1.7520 0.9400 ;
      RECT 1.1700 0.5710 1.9560 0.6210 ;
      RECT 1.7020 0.6210 1.7520 0.8900 ;
      RECT 1.1130 0.9400 1.1630 1.0080 ;
      RECT 0.8710 1.0080 1.1630 1.0580 ;
      RECT 1.1700 0.4580 1.2200 0.5710 ;
      RECT 0.8710 0.4080 1.2200 0.4580 ;
      RECT 1.7990 1.1580 1.8490 1.3200 ;
      RECT 0.4310 1.1080 1.8490 1.1580 ;
      RECT 0.4310 1.1580 0.4810 1.3200 ;
      RECT 0.4310 0.1530 1.2410 0.2030 ;
      RECT 1.1910 0.2030 1.2410 0.3260 ;
      RECT 0.4310 0.2030 0.4810 0.3260 ;
      RECT 1.4640 0.3710 1.8800 0.4210 ;
    LAYER PO ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 1.2770 0.0680 1.3070 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
  END
END XOR2X2_LVT

MACRO XOR3X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.256 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.2560 1.7020 ;
        RECT 0.7350 1.2180 0.7850 1.6420 ;
        RECT 1.9510 1.2180 2.0010 1.6420 ;
        RECT 1.1910 1.2180 1.2410 1.6420 ;
        RECT 0.4310 1.2230 0.4810 1.6420 ;
        RECT 2.7110 1.2150 2.7610 1.6420 ;
        RECT 3.7750 1.4070 3.8250 1.6420 ;
        RECT 3.4550 1.3570 3.8250 1.4070 ;
    END
  END VDD

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.5460 0.8570 3.7050 0.9730 ;
        RECT 3.5470 0.6690 3.5970 0.8570 ;
        RECT 3.0910 0.6190 3.5970 0.6690 ;
        RECT 3.0910 0.6690 3.1410 0.7310 ;
    END
    ANTENNAGATEAREA 0.0498 ;
  END A3

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.9270 1.2490 4.0570 1.2990 ;
        RECT 3.9270 1.2990 3.9770 1.5460 ;
        RECT 4.0070 1.1190 4.0570 1.2490 ;
        RECT 4.0070 1.0090 4.1590 1.1190 ;
        RECT 4.0070 0.5420 4.0570 1.0090 ;
        RECT 3.9270 0.4920 4.0570 0.5420 ;
        RECT 3.9270 0.1270 3.9770 0.4920 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.2560 0.0300 ;
        RECT 2.7110 0.0300 2.7610 0.3260 ;
        RECT 2.1910 0.0300 2.2410 0.2630 ;
        RECT 0.1620 0.0300 0.2120 0.3910 ;
        RECT 3.7750 0.0300 3.8250 0.2110 ;
        RECT 1.9200 0.2630 2.2410 0.3130 ;
        RECT 0.1620 0.3910 0.7330 0.4410 ;
        RECT 3.4500 0.2110 3.8430 0.2610 ;
        RECT 0.4310 0.3000 0.4810 0.3910 ;
        RECT 0.6830 0.3200 0.7330 0.3910 ;
        RECT 0.6830 0.2700 1.2720 0.3200 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1140 0.6640 1.7720 0.7140 ;
        RECT 1.1140 0.5530 1.2710 0.6640 ;
        RECT 1.7220 0.6420 1.7720 0.6640 ;
        RECT 1.7220 0.5920 2.5330 0.6420 ;
        RECT 2.4830 0.6420 2.5330 0.7540 ;
    END
    ANTENNAGATEAREA 0.0783 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8120 0.7050 0.9670 0.8030 ;
        RECT 0.8120 0.8030 2.0770 0.8530 ;
        RECT 2.0270 0.7030 2.0770 0.8030 ;
        RECT 1.8750 0.7030 1.9250 0.8030 ;
    END
    ANTENNAGATEAREA 0.0753 ;
  END A2
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 4.3710 1.7730 ;
    LAYER M1 ;
      RECT 3.3210 1.5340 3.4610 1.5840 ;
      RECT 2.5590 1.1650 2.6090 1.3050 ;
      RECT 2.5590 1.0580 2.6090 1.1150 ;
      RECT 1.4640 1.0080 2.6090 1.0580 ;
      RECT 2.5590 0.8590 2.6090 1.0080 ;
      RECT 2.5590 0.2410 2.6090 0.4640 ;
      RECT 3.3210 1.2990 3.3710 1.5340 ;
      RECT 3.0070 1.2490 3.3850 1.2990 ;
      RECT 3.0070 1.1650 3.0570 1.2490 ;
      RECT 2.5590 1.1150 3.0570 1.1650 ;
      RECT 2.5590 0.8090 2.6640 0.8590 ;
      RECT 2.6140 0.6540 2.6640 0.8090 ;
      RECT 2.6140 0.6040 2.8370 0.6540 ;
      RECT 2.6140 0.5140 2.6640 0.6040 ;
      RECT 2.7870 0.6540 2.8370 0.6850 ;
      RECT 2.7870 0.5730 2.8370 0.6040 ;
      RECT 1.5300 0.4640 2.6640 0.5140 ;
      RECT 1.5300 0.3750 1.5800 0.4640 ;
      RECT 1.4790 0.3250 1.5800 0.3750 ;
      RECT 0.3970 1.0180 0.9530 1.0680 ;
      RECT 0.8870 0.3770 0.9370 0.4910 ;
      RECT 0.3970 0.4910 0.9370 0.5410 ;
      RECT 0.3970 0.6540 0.4470 1.0180 ;
      RECT 0.3390 0.6040 0.5730 0.6540 ;
      RECT 0.3970 0.5410 0.4470 0.6040 ;
      RECT 0.9990 0.4080 1.4080 0.4580 ;
      RECT 1.3580 0.4580 1.4080 0.5640 ;
      RECT 0.6320 0.9180 1.0890 0.9680 ;
      RECT 1.0390 0.9680 1.0890 1.0680 ;
      RECT 1.3580 0.5640 1.6540 0.6140 ;
      RECT 0.9990 0.4580 1.0490 0.5910 ;
      RECT 0.6320 0.5910 1.0490 0.6410 ;
      RECT 0.6320 0.6410 0.6820 0.9180 ;
      RECT 0.2790 0.1530 1.6970 0.2030 ;
      RECT 1.3430 0.2030 1.3930 0.3000 ;
      RECT 1.6470 0.2030 1.6970 0.3000 ;
      RECT 0.5830 0.2030 0.6330 0.3410 ;
      RECT 0.2790 0.2030 0.3290 0.3410 ;
      RECT 3.5920 0.4180 3.7450 0.4680 ;
      RECT 3.6950 0.4680 3.7450 0.7100 ;
      RECT 3.6950 0.7100 3.8220 0.7600 ;
      RECT 3.7720 0.7600 3.8220 1.0290 ;
      RECT 3.2980 1.0290 3.8220 1.0790 ;
      RECT 3.2980 0.7690 3.3480 1.0290 ;
      RECT 3.2120 0.7190 3.3480 0.7690 ;
      RECT 1.7830 0.3640 2.4880 0.4140 ;
      RECT 3.8210 0.6040 3.9320 0.6540 ;
      RECT 3.8810 0.6540 3.9310 1.1490 ;
      RECT 3.1500 1.1490 3.9310 1.1990 ;
      RECT 2.9870 0.5690 3.0370 0.8220 ;
      RECT 3.1800 0.8720 3.2300 1.1490 ;
      RECT 2.9870 0.8220 3.2300 0.8720 ;
      RECT 3.4350 0.3680 3.4850 0.5190 ;
      RECT 3.1310 0.3180 3.4850 0.3680 ;
      RECT 2.9870 0.5190 3.4850 0.5690 ;
      RECT 2.4070 1.1680 2.4570 1.3200 ;
      RECT 0.2790 1.1180 2.4570 1.1680 ;
      RECT 0.2790 1.1680 0.3290 1.3200 ;
      RECT 0.5830 1.1680 0.6330 1.3200 ;
      RECT 3.0150 0.1110 3.4610 0.1610 ;
      RECT 3.0150 0.1610 3.0650 0.3260 ;
      RECT 2.8270 0.9800 3.0960 1.0300 ;
      RECT 2.8470 0.4180 3.3850 0.4680 ;
      RECT 2.8870 0.4680 2.9370 0.9800 ;
      RECT 1.3270 0.9040 2.1690 0.9540 ;
    LAYER PO ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 3.7090 0.0680 3.7390 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 1.2770 0.0680 1.3070 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
  END
END XOR3X1_LVT

MACRO XOR3X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.408 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.9270 0.9670 3.9770 1.5460 ;
        RECT 3.9270 0.9170 4.1930 0.9670 ;
        RECT 4.0490 0.8560 4.1930 0.9170 ;
        RECT 4.1430 0.4950 4.1930 0.8560 ;
        RECT 3.9270 0.4450 4.1930 0.4950 ;
        RECT 3.9270 0.1280 3.9770 0.4450 ;
    END
    ANTENNADIFFAREA 0.1464 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0260 0.6270 2.0760 0.7050 ;
        RECT 2.0260 0.7050 2.1830 0.8290 ;
        RECT 2.0260 0.5770 2.5640 0.6270 ;
    END
    ANTENNAGATEAREA 0.0765 ;
  END A1

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4410 1.5110 3.5980 1.5750 ;
        RECT 3.0600 1.4610 3.5990 1.5110 ;
    END
    ANTENNAGATEAREA 0.036 ;
  END A3

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.4080 1.7020 ;
        RECT 4.0790 1.3560 4.1290 1.6420 ;
        RECT 2.7110 1.0830 2.7610 1.6420 ;
        RECT 0.4310 1.2600 0.4810 1.6420 ;
        RECT 0.8870 1.2180 0.9370 1.6420 ;
        RECT 2.1080 1.2560 2.1580 1.6420 ;
        RECT 3.7750 1.1410 3.8250 1.6420 ;
        RECT 1.6110 1.2060 2.1690 1.2560 ;
        RECT 3.4550 1.0910 3.8250 1.1410 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.4080 0.0300 ;
        RECT 3.7750 0.0300 3.8250 0.2000 ;
        RECT 4.0790 0.0300 4.1290 0.2250 ;
        RECT 2.7110 0.0300 2.7610 0.0910 ;
        RECT 0.1350 0.0300 0.1850 0.3120 ;
        RECT 2.7110 0.0910 3.4760 0.1410 ;
        RECT 0.1350 0.3120 0.9760 0.3620 ;
        RECT 2.7110 0.1410 2.7610 0.2660 ;
        RECT 0.9260 0.3620 0.9760 0.4450 ;
        RECT 0.9260 0.4450 1.5130 0.4950 ;
        RECT 1.4630 0.3620 1.5130 0.4450 ;
        RECT 1.4630 0.3120 2.1840 0.3620 ;
    END
  END VSS

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8100 0.5530 0.9670 0.6630 ;
        RECT 0.8100 0.6630 0.8600 0.7320 ;
        RECT 0.8100 0.7320 1.7970 0.7820 ;
    END
    ANTENNAGATEAREA 0.0735 ;
  END A2
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 4.5230 1.7810 ;
    LAYER M1 ;
      RECT 2.5590 0.4530 2.6660 0.5030 ;
      RECT 2.6160 0.5030 2.6660 0.6480 ;
      RECT 2.6160 0.6480 2.8780 0.6980 ;
      RECT 2.6160 0.6980 2.6660 0.8630 ;
      RECT 2.5590 0.8630 2.6660 0.9130 ;
      RECT 2.5590 0.9830 3.3850 1.0060 ;
      RECT 1.4190 1.0060 3.3850 1.0330 ;
      RECT 2.2390 0.3160 3.0840 0.3660 ;
      RECT 1.1910 0.1530 1.2410 0.2350 ;
      RECT 1.4190 0.9340 1.4690 1.0060 ;
      RECT 1.1550 0.8840 1.4690 0.9340 ;
      RECT 2.5590 0.3660 2.6090 0.4530 ;
      RECT 2.5590 0.1530 2.6090 0.3160 ;
      RECT 1.1910 0.1030 2.6090 0.1530 ;
      RECT 2.5590 0.9130 2.6090 0.9830 ;
      RECT 1.4190 1.0330 2.6090 1.0560 ;
      RECT 2.5590 1.0560 2.6090 1.2640 ;
      RECT 0.2530 0.1960 1.0890 0.2460 ;
      RECT 1.0390 0.1630 1.0890 0.1960 ;
      RECT 1.0390 0.2460 1.0890 0.3340 ;
      RECT 1.0390 0.3340 1.3930 0.3840 ;
      RECT 1.3430 0.2460 1.3930 0.3340 ;
      RECT 1.8910 0.4120 2.0370 0.4620 ;
      RECT 1.8910 0.9060 2.0350 0.9560 ;
      RECT 1.8910 0.4620 1.9410 0.6050 ;
      RECT 1.0830 0.6050 1.9410 0.6550 ;
      RECT 1.8910 0.6550 1.9410 0.9060 ;
      RECT 2.8270 0.8830 3.0810 0.9330 ;
      RECT 2.9360 0.4660 2.9860 0.8830 ;
      RECT 2.8270 0.4160 3.4000 0.4660 ;
      RECT 1.0390 1.4480 1.8660 1.4980 ;
      RECT 1.0390 1.2180 1.0890 1.4480 ;
      RECT 1.3430 1.2180 1.3930 1.4480 ;
      RECT 1.4950 1.2170 1.5450 1.4480 ;
      RECT 3.2430 0.7430 3.7250 0.7930 ;
      RECT 3.2430 0.6490 3.2930 0.7430 ;
      RECT 3.6230 0.7930 3.6730 0.9320 ;
      RECT 3.6750 0.4690 3.7250 0.7430 ;
      RECT 3.5920 0.4190 3.7250 0.4690 ;
      RECT 3.7850 0.6040 4.0840 0.6540 ;
      RECT 3.7850 0.6540 3.8350 0.9910 ;
      RECT 3.7850 0.3560 3.8350 0.6040 ;
      RECT 3.4900 0.9910 3.8350 1.0410 ;
      RECT 3.1490 0.3060 3.8350 0.3560 ;
      RECT 3.4900 0.9270 3.5400 0.9910 ;
      RECT 3.1460 0.8770 3.5400 0.9270 ;
      RECT 3.4710 0.4190 3.5210 0.5770 ;
      RECT 3.3790 0.5770 3.5210 0.6270 ;
      RECT 2.4070 1.1560 2.4570 1.2670 ;
      RECT 0.2790 1.1060 2.4570 1.1560 ;
      RECT 0.2790 1.1560 0.3290 1.4610 ;
      RECT 0.5830 1.1560 0.6330 1.4610 ;
      RECT 0.6530 0.9700 0.8160 1.0200 ;
      RECT 0.6530 0.4240 0.8160 0.4740 ;
      RECT 0.6530 0.6540 0.7030 0.9700 ;
      RECT 0.3240 0.6040 0.7030 0.6540 ;
      RECT 0.6530 0.4740 0.7030 0.6040 ;
      RECT 1.4790 0.2070 2.4880 0.2570 ;
    LAYER PO ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 1.2770 0.0680 1.3070 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 3.7090 0.0680 3.7390 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 4.3170 0.0680 4.3470 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
  END
END XOR3X2_LVT

MACRO SDFFSSRX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.472 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 5.4720 1.7020 ;
        RECT 4.9910 0.9470 5.0410 1.6420 ;
        RECT 2.1030 1.3520 2.1530 1.6420 ;
        RECT 4.7270 1.4660 4.7770 1.6420 ;
        RECT 1.1510 1.2850 1.2010 1.6420 ;
        RECT 0.2790 1.3460 0.3290 1.6420 ;
        RECT 3.4710 1.3660 3.5210 1.6420 ;
        RECT 2.1030 1.3020 2.4730 1.3520 ;
        RECT 4.2150 1.4160 4.7770 1.4660 ;
        RECT 1.1510 1.2350 1.2570 1.2850 ;
        RECT 0.2790 1.2960 0.6330 1.3460 ;
        RECT 3.3190 1.3160 3.5210 1.3660 ;
        RECT 4.6870 1.1920 4.7370 1.4160 ;
        RECT 0.2790 0.9300 0.3290 1.2960 ;
        RECT 0.5830 0.9800 0.6330 1.2960 ;
        RECT 3.3190 1.1520 3.3690 1.3160 ;
    END
  END VDD

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.1130 0.4270 5.2230 0.5110 ;
        RECT 4.8390 0.3770 5.2230 0.4270 ;
        RECT 5.1730 0.5110 5.2230 0.8080 ;
        RECT 4.8390 0.1360 4.8890 0.3770 ;
        RECT 4.8390 0.8080 5.2230 0.8580 ;
        RECT 4.8390 0.8580 4.8890 1.5460 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.1430 1.0690 5.3750 1.1190 ;
        RECT 5.2650 1.0090 5.3750 1.0690 ;
        RECT 5.1430 1.1190 5.1930 1.5460 ;
        RECT 5.3250 0.3100 5.3750 1.0090 ;
        RECT 5.1430 0.2600 5.3750 0.3100 ;
        RECT 5.1430 0.1360 5.1930 0.2600 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7010 0.4210 0.7510 ;
        RECT 0.2490 0.7510 0.3590 0.8250 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SETB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2250 1.4650 2.3970 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 5.4720 0.0300 ;
        RECT 4.1910 0.0300 4.2410 0.2040 ;
        RECT 0.2790 0.0300 0.3290 0.3550 ;
        RECT 2.0630 0.0300 2.1130 0.3010 ;
        RECT 1.1910 0.0300 1.2410 0.3590 ;
        RECT 4.9910 0.0300 5.0410 0.3030 ;
        RECT 4.6870 0.0300 4.7370 0.4010 ;
        RECT 4.1910 0.2040 4.2970 0.2540 ;
        RECT 0.2790 0.3550 0.6330 0.4050 ;
        RECT 2.0630 0.3010 3.5210 0.3510 ;
        RECT 0.5830 0.4050 0.6330 0.5290 ;
        RECT 0.2790 0.4050 0.3290 0.5130 ;
        RECT 3.4710 0.3510 3.5210 0.4750 ;
        RECT 2.4070 0.3510 2.4570 0.5760 ;
        RECT 3.3190 0.3510 3.3690 0.4750 ;
    END
  END VSS

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0290 0.8280 2.1830 0.9670 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9470 0.5530 1.1190 0.6730 ;
    END
    ANTENNAGATEAREA 0.0255 ;
  END D

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2510 1.4160 1.6370 1.4660 ;
        RECT 1.3130 1.3130 1.4230 1.4160 ;
    END
    ANTENNAGATEAREA 0.039 ;
  END SE

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 0.0970 0.5110 0.2010 ;
        RECT 0.4010 0.2010 0.7250 0.2510 ;
    END
    ANTENNAGATEAREA 0.0255 ;
  END RSTB
  OBS
    LAYER PO ;
      RECT 0.2130 0.0760 0.2430 1.6060 ;
      RECT 0.3650 0.0760 0.3950 1.6060 ;
      RECT 3.2530 0.9660 3.2830 1.6060 ;
      RECT 2.3410 0.0760 2.3710 1.6060 ;
      RECT 5.3810 0.0760 5.4110 1.6060 ;
      RECT 3.4050 0.0760 3.4350 1.6060 ;
      RECT 1.7330 0.0760 1.7630 0.6000 ;
      RECT 0.8210 0.8380 0.8510 1.6060 ;
      RECT 1.1250 0.0760 1.1550 1.6060 ;
      RECT 2.7970 0.0760 2.8270 0.5970 ;
      RECT 3.8610 1.0320 3.8910 1.6060 ;
      RECT 5.2290 0.0760 5.2590 1.6060 ;
      RECT 0.5170 0.0760 0.5470 1.6060 ;
      RECT 1.5810 0.8700 1.6110 1.6060 ;
      RECT 4.6210 0.0760 4.6510 0.7550 ;
      RECT 4.7730 0.0760 4.8030 1.6060 ;
      RECT 0.8210 0.0760 0.8510 0.6510 ;
      RECT 2.7970 0.9200 2.8270 1.6060 ;
      RECT 2.6450 0.0760 2.6750 1.6060 ;
      RECT 0.0610 0.0760 0.0910 1.6060 ;
      RECT 1.5810 0.0760 1.6110 0.6000 ;
      RECT 3.1010 0.0760 3.1310 1.6060 ;
      RECT 1.2770 0.0760 1.3070 1.6060 ;
      RECT 1.4290 0.0760 1.4590 1.6060 ;
      RECT 1.8850 0.0760 1.9150 1.6060 ;
      RECT 4.9250 0.0760 4.9550 1.6060 ;
      RECT 2.4930 0.0760 2.5230 1.6060 ;
      RECT 3.5570 0.0760 3.5870 1.6060 ;
      RECT 4.6210 1.1320 4.6510 1.6060 ;
      RECT 3.2530 0.0760 3.2830 0.7510 ;
      RECT 4.1650 0.0760 4.1950 1.6060 ;
      RECT 4.4690 0.0760 4.4990 1.6060 ;
      RECT 2.9490 0.0760 2.9790 1.6060 ;
      RECT 5.0770 0.0760 5.1070 1.6060 ;
      RECT 4.3170 0.0760 4.3470 1.6060 ;
      RECT 2.1890 0.0760 2.2190 1.6060 ;
      RECT 3.8610 0.0760 3.8910 0.5970 ;
      RECT 3.7090 0.0760 3.7390 1.6060 ;
      RECT 0.6690 0.0760 0.6990 0.5970 ;
      RECT 0.6690 0.8160 0.6990 1.6060 ;
      RECT 4.0130 0.0760 4.0430 1.6060 ;
      RECT 0.9730 0.0760 1.0030 1.6060 ;
      RECT 2.0370 0.0760 2.0670 1.6060 ;
      RECT 1.7330 0.8700 1.7630 1.6060 ;
    LAYER NWELL ;
      RECT -0.1150 0.6790 5.5870 1.7730 ;
    LAYER M1 ;
      RECT 4.3920 0.1540 4.4420 0.3040 ;
      RECT 4.0390 0.3040 4.4420 0.3540 ;
      RECT 4.2910 0.1040 4.5250 0.1540 ;
      RECT 4.0390 0.3540 4.0890 0.8080 ;
      RECT 4.0390 0.8080 4.1290 0.8580 ;
      RECT 4.0790 0.8580 4.1290 1.1660 ;
      RECT 2.7110 0.7260 2.8010 0.7760 ;
      RECT 2.7110 0.7760 2.7610 1.2020 ;
      RECT 2.7510 0.5760 2.8010 0.7260 ;
      RECT 1.6470 1.2020 2.7610 1.2520 ;
      RECT 2.7110 0.5260 2.8010 0.5760 ;
      RECT 2.7110 0.4300 2.7610 0.5260 ;
      RECT 1.6470 0.3490 1.6970 1.2020 ;
      RECT 2.9630 0.6730 3.3090 0.7230 ;
      RECT 2.9630 0.8800 3.1650 0.9300 ;
      RECT 2.9630 0.7230 3.0130 0.8800 ;
      RECT 3.1150 0.9300 3.1650 1.3170 ;
      RECT 2.8230 1.3170 3.1650 1.3670 ;
      RECT 2.8230 1.3670 2.8730 1.5280 ;
      RECT 2.6190 1.5280 2.8730 1.5780 ;
      RECT 2.1630 0.6260 2.5490 0.6760 ;
      RECT 2.2550 0.6760 2.3050 1.1520 ;
      RECT 2.2550 0.4010 2.3050 0.6260 ;
      RECT 1.7990 1.1020 2.0170 1.1520 ;
      RECT 1.7990 0.3490 2.0010 0.3990 ;
      RECT 1.9510 0.3990 2.0010 0.5370 ;
      RECT 1.7990 0.3990 1.8490 1.1020 ;
      RECT 3.9210 0.1040 4.0690 0.1510 ;
      RECT 3.2270 0.1510 4.0690 0.1540 ;
      RECT 3.2270 0.1540 3.9710 0.2010 ;
      RECT 0.7000 0.5730 0.8770 0.6230 ;
      RECT 0.7000 0.6230 0.7500 0.8120 ;
      RECT 0.4310 0.8120 0.7500 0.8620 ;
      RECT 0.4310 0.8620 0.4810 1.2460 ;
      RECT 0.4310 0.4550 0.4810 0.6010 ;
      RECT 0.4710 0.6510 0.5210 0.8120 ;
      RECT 0.4310 0.6010 0.5210 0.6510 ;
      RECT 4.5870 0.6770 4.6770 0.7270 ;
      RECT 4.5870 0.7270 4.6370 1.3160 ;
      RECT 3.8750 1.3160 4.6370 1.3660 ;
      RECT 3.8750 1.3660 3.9250 1.5280 ;
      RECT 3.6310 1.5280 3.9250 1.5780 ;
      RECT 3.6310 1.2660 3.6810 1.5280 ;
      RECT 3.4670 1.0440 3.5170 1.2160 ;
      RECT 3.2270 0.9940 3.5170 1.0440 ;
      RECT 3.4670 1.2160 3.6810 1.2660 ;
      RECT 4.8150 0.7080 5.1170 0.7580 ;
      RECT 5.0670 0.6210 5.1170 0.7080 ;
      RECT 4.8150 0.6270 4.8650 0.7080 ;
      RECT 4.4430 0.5770 4.8650 0.6270 ;
      RECT 3.9870 1.5280 4.6770 1.5780 ;
      RECT 1.2910 0.3190 1.3930 0.3690 ;
      RECT 1.3430 0.3690 1.3930 1.0020 ;
      RECT 1.2910 0.1510 1.3410 0.3190 ;
      RECT 1.2910 0.1010 1.9410 0.1510 ;
      RECT 0.7190 0.3010 1.1050 0.3510 ;
      RECT 0.8710 0.4430 1.2500 0.4930 ;
      RECT 1.2000 0.4930 1.2500 1.0520 ;
      RECT 0.8870 1.0520 1.5450 1.1020 ;
      RECT 1.4950 1.1020 1.5450 1.2520 ;
      RECT 1.4950 0.3490 1.5450 1.0520 ;
      RECT 0.8870 1.1020 0.9370 1.2460 ;
      RECT 0.8870 0.9800 0.9370 1.0520 ;
      RECT 1.4030 0.2040 1.7890 0.2540 ;
      RECT 0.7350 1.3160 1.0890 1.3660 ;
      RECT 0.7350 0.9800 0.7850 1.3160 ;
      RECT 1.0390 1.1920 1.0890 1.3160 ;
      RECT 1.7070 1.4160 1.9460 1.4660 ;
      RECT 2.1630 0.1040 3.0050 0.1540 ;
      RECT 2.7870 0.1540 2.8370 0.2170 ;
      RECT 2.9230 1.4170 3.3090 1.4670 ;
      RECT 2.5590 0.7260 2.6610 0.7760 ;
      RECT 2.5590 0.7760 2.6090 1.1520 ;
      RECT 2.6110 0.6760 2.6610 0.7260 ;
      RECT 2.6110 0.6260 2.7010 0.6760 ;
      RECT 2.6110 0.4960 2.6610 0.6260 ;
      RECT 2.5430 0.4460 2.6610 0.4960 ;
      RECT 4.9150 0.5270 4.9650 0.6580 ;
      RECT 4.3430 0.4770 4.9650 0.5270 ;
      RECT 3.9270 0.3000 3.9770 1.2160 ;
      RECT 4.3430 0.5270 4.3930 0.6540 ;
      RECT 4.1390 0.6540 4.3930 0.6770 ;
      RECT 4.1390 0.6770 4.4730 0.7040 ;
      RECT 4.3430 0.7040 4.4730 0.7270 ;
      RECT 4.4230 0.7270 4.4730 1.2160 ;
      RECT 3.9270 1.2160 4.4730 1.2660 ;
      RECT 2.8630 0.5730 3.6130 0.6230 ;
      RECT 3.0150 0.4300 3.0650 0.5730 ;
      RECT 2.8630 0.6230 2.9130 1.1960 ;
      RECT 2.8630 0.4300 2.9130 0.5730 ;
      RECT 2.8630 1.1960 3.0650 1.2460 ;
      RECT 3.0150 1.1380 3.0650 1.1960 ;
      RECT 0.4910 1.5340 0.8770 1.5840 ;
      RECT 3.0700 0.7730 3.8250 0.8230 ;
      RECT 3.6230 0.8230 3.6730 1.1660 ;
      RECT 3.7750 0.8230 3.8250 1.3800 ;
      RECT 3.7750 0.5020 3.8250 0.7730 ;
      RECT 3.6230 0.4520 3.8250 0.5020 ;
      RECT 3.6230 0.3000 3.6730 0.4520 ;
      RECT 3.7750 0.3000 3.8250 0.4520 ;
  END
END SDFFSSRX1_LVT

MACRO SDFFSSRX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.776 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 5.7760 1.7020 ;
        RECT 5.1430 0.9600 5.1930 1.6420 ;
        RECT 4.8390 0.9120 4.8890 1.6420 ;
        RECT 5.4470 1.0520 5.4970 1.6420 ;
        RECT 2.1030 1.3520 2.1530 1.6420 ;
        RECT 4.7270 1.4660 4.7770 1.6420 ;
        RECT 1.1510 1.2850 1.2010 1.6420 ;
        RECT 0.2790 1.3460 0.3290 1.6420 ;
        RECT 3.4710 1.3660 3.5210 1.6420 ;
        RECT 2.1030 1.3020 2.4730 1.3520 ;
        RECT 4.2150 1.4160 4.7770 1.4660 ;
        RECT 1.1510 1.2350 1.2570 1.2850 ;
        RECT 0.2790 1.2960 0.6330 1.3460 ;
        RECT 3.3190 1.3160 3.5210 1.3660 ;
        RECT 4.6870 1.1920 4.7370 1.4160 ;
        RECT 0.2790 0.9300 0.3290 1.2960 ;
        RECT 0.5830 0.9800 0.6330 1.2960 ;
        RECT 3.3190 1.1730 3.3690 1.3160 ;
    END
  END VDD

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7010 0.4210 0.7510 ;
        RECT 0.2490 0.7510 0.3590 0.8250 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SETB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2250 1.4650 2.3970 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 5.7760 0.0300 ;
        RECT 4.1910 0.0300 4.2410 0.2040 ;
        RECT 0.2790 0.0300 0.3290 0.3550 ;
        RECT 2.0630 0.0300 2.1130 0.3010 ;
        RECT 1.1910 0.0300 1.2410 0.3590 ;
        RECT 4.6870 0.0300 4.7370 0.4010 ;
        RECT 5.4470 0.0300 5.4970 0.2200 ;
        RECT 5.1430 0.0300 5.1930 0.3190 ;
        RECT 4.8390 0.0300 4.8890 0.4080 ;
        RECT 4.1910 0.2040 4.2970 0.2540 ;
        RECT 0.2790 0.3550 0.6330 0.4050 ;
        RECT 2.0630 0.3010 3.5210 0.3510 ;
        RECT 0.5830 0.4050 0.6330 0.5290 ;
        RECT 0.2790 0.4050 0.3290 0.5130 ;
        RECT 3.4710 0.3510 3.5210 0.4750 ;
        RECT 2.4070 0.3510 2.4570 0.5760 ;
        RECT 3.3190 0.3510 3.3690 0.4750 ;
    END
  END VSS

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0290 0.8280 2.1830 0.9670 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9470 0.5530 1.1190 0.6730 ;
    END
    ANTENNAGATEAREA 0.0255 ;
  END D

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2510 1.4160 1.6370 1.4660 ;
        RECT 1.3130 1.3130 1.4230 1.4160 ;
    END
    ANTENNAGATEAREA 0.039 ;
  END SE

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.5690 0.0970 5.6790 0.2070 ;
        RECT 5.6110 0.2070 5.6610 0.2700 ;
        RECT 5.2950 0.2700 5.6610 0.3200 ;
        RECT 5.2950 0.1480 5.3450 0.2700 ;
        RECT 5.6110 0.3200 5.6610 0.9180 ;
        RECT 5.2950 0.9180 5.6610 0.9680 ;
        RECT 5.2950 0.9680 5.3450 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 0.0970 0.5110 0.2010 ;
        RECT 0.4010 0.2010 0.7250 0.2510 ;
    END
    ANTENNAGATEAREA 0.0255 ;
  END RSTB

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.9910 0.1480 5.0410 0.3740 ;
        RECT 4.9910 0.3740 5.5370 0.4240 ;
        RECT 5.4170 0.4240 5.5370 0.5110 ;
        RECT 5.4870 0.5110 5.5370 0.8040 ;
        RECT 4.9910 0.8040 5.5370 0.8540 ;
        RECT 4.9910 0.8540 5.0410 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q
  OBS
    LAYER PO ;
      RECT 2.9490 0.0760 2.9790 1.6060 ;
      RECT 4.3170 0.0760 4.3470 1.6060 ;
      RECT 2.1890 0.0760 2.2190 1.6060 ;
      RECT 3.8610 0.0760 3.8910 0.5970 ;
      RECT 3.7090 0.0760 3.7390 1.6060 ;
      RECT 0.6690 0.0760 0.6990 0.5970 ;
      RECT 0.6690 0.8020 0.6990 1.6060 ;
      RECT 4.0130 0.0760 4.0430 1.6060 ;
      RECT 0.9730 0.0760 1.0030 1.6060 ;
      RECT 2.0370 0.0760 2.0670 1.6060 ;
      RECT 1.7330 0.8700 1.7630 1.6060 ;
      RECT 5.5330 0.0680 5.5630 1.6060 ;
      RECT 0.2130 0.0760 0.2430 1.6060 ;
      RECT 0.3650 0.0760 0.3950 1.6060 ;
      RECT 3.2530 0.9660 3.2830 1.6060 ;
      RECT 2.3410 0.0760 2.3710 1.6060 ;
      RECT 3.4050 0.0760 3.4350 1.6060 ;
      RECT 1.7330 0.0760 1.7630 0.6000 ;
      RECT 0.8210 0.8340 0.8510 1.6060 ;
      RECT 1.1250 0.0760 1.1550 1.6060 ;
      RECT 4.7730 0.0680 4.8030 1.6060 ;
      RECT 2.7970 0.0760 2.8270 0.5970 ;
      RECT 3.8610 1.0320 3.8910 1.6060 ;
      RECT 0.5170 0.0760 0.5470 1.6060 ;
      RECT 1.5810 0.8700 1.6110 1.6060 ;
      RECT 4.6210 0.0760 4.6510 0.7550 ;
      RECT 5.6850 0.0680 5.7150 1.6060 ;
      RECT 0.8210 0.0760 0.8510 0.6510 ;
      RECT 2.7970 0.9200 2.8270 1.6060 ;
      RECT 2.6450 0.0760 2.6750 1.6060 ;
      RECT 4.9250 0.0680 4.9550 1.6060 ;
      RECT 5.2290 0.0680 5.2590 1.6060 ;
      RECT 0.0610 0.0760 0.0910 1.6060 ;
      RECT 1.5810 0.0760 1.6110 0.6000 ;
      RECT 5.3810 0.0680 5.4110 1.6060 ;
      RECT 5.0770 0.0680 5.1070 1.6060 ;
      RECT 3.1010 0.0760 3.1310 1.6060 ;
      RECT 1.2770 0.0760 1.3070 1.6060 ;
      RECT 1.4290 0.0760 1.4590 1.6060 ;
      RECT 1.8850 0.0760 1.9150 1.6060 ;
      RECT 2.4930 0.0760 2.5230 1.6060 ;
      RECT 3.5570 0.0760 3.5870 1.6060 ;
      RECT 4.6210 1.1320 4.6510 1.6060 ;
      RECT 3.2530 0.0760 3.2830 0.7510 ;
      RECT 4.1650 0.0760 4.1950 1.6060 ;
      RECT 4.4690 0.0760 4.4990 1.6060 ;
    LAYER NWELL ;
      RECT -0.1150 0.6790 5.8910 1.7730 ;
    LAYER M1 ;
      RECT 4.3920 0.1540 4.4420 0.3040 ;
      RECT 4.0390 0.3040 4.4420 0.3540 ;
      RECT 4.2910 0.1040 4.5250 0.1540 ;
      RECT 4.0390 0.3540 4.0890 0.8080 ;
      RECT 4.0390 0.8080 4.1290 0.8580 ;
      RECT 4.0790 0.8580 4.1290 1.1660 ;
      RECT 2.9630 0.6730 3.3090 0.7230 ;
      RECT 2.9630 0.8800 3.1650 0.9300 ;
      RECT 3.1150 0.9300 3.1650 1.3170 ;
      RECT 2.9630 0.7230 3.0130 0.8800 ;
      RECT 2.8230 1.3170 3.1650 1.3670 ;
      RECT 2.8230 1.3670 2.8730 1.5280 ;
      RECT 2.6190 1.5280 2.8730 1.5780 ;
      RECT 3.0700 0.7730 3.8250 0.8230 ;
      RECT 3.6230 0.8230 3.6730 1.1660 ;
      RECT 3.7750 0.8230 3.8250 1.3800 ;
      RECT 3.7750 0.5020 3.8250 0.7730 ;
      RECT 3.6230 0.4520 3.8250 0.5020 ;
      RECT 3.7750 0.3000 3.8250 0.4520 ;
      RECT 3.6230 0.3000 3.6730 0.4520 ;
      RECT 0.8870 1.0520 1.5450 1.1020 ;
      RECT 1.4950 1.1020 1.5450 1.2520 ;
      RECT 1.4950 0.3490 1.5450 1.0520 ;
      RECT 1.2000 0.4930 1.2500 1.0520 ;
      RECT 0.8710 0.4430 1.2500 0.4930 ;
      RECT 0.8870 1.1020 0.9370 1.2460 ;
      RECT 0.8870 0.9800 0.9370 1.0520 ;
      RECT 3.2270 0.1540 3.9710 0.2010 ;
      RECT 3.2270 0.1510 4.0690 0.1540 ;
      RECT 3.9210 0.1040 4.0690 0.1510 ;
      RECT 4.5870 0.6770 4.6770 0.7270 ;
      RECT 4.5870 0.7270 4.6370 1.3160 ;
      RECT 3.8750 1.3160 4.6370 1.3660 ;
      RECT 3.8750 1.3660 3.9250 1.5280 ;
      RECT 3.6310 1.5280 3.9250 1.5780 ;
      RECT 3.6310 1.2660 3.6810 1.5280 ;
      RECT 3.4670 1.0440 3.5170 1.2160 ;
      RECT 3.2270 0.9940 3.5170 1.0440 ;
      RECT 3.4670 1.2160 3.6810 1.2660 ;
      RECT 2.8630 0.5730 3.6130 0.6230 ;
      RECT 3.0150 0.4300 3.0650 0.5730 ;
      RECT 2.8630 0.6230 2.9130 1.1960 ;
      RECT 2.8630 0.4300 2.9130 0.5730 ;
      RECT 2.8630 1.1960 3.0650 1.2460 ;
      RECT 3.0150 1.1420 3.0650 1.1960 ;
      RECT 0.4910 1.5340 0.8770 1.5840 ;
      RECT 2.7110 0.7260 2.8010 0.7760 ;
      RECT 2.7110 0.7760 2.7610 1.2020 ;
      RECT 2.7510 0.5760 2.8010 0.7260 ;
      RECT 1.6470 1.2020 2.7610 1.2520 ;
      RECT 2.7110 0.5260 2.8010 0.5760 ;
      RECT 2.7110 0.4300 2.7610 0.5260 ;
      RECT 1.6470 0.3490 1.6970 1.2020 ;
      RECT 2.1630 0.6260 2.5490 0.6760 ;
      RECT 2.2550 0.6760 2.3050 1.1520 ;
      RECT 2.2550 0.4010 2.3050 0.6260 ;
      RECT 1.7990 1.1020 2.0170 1.1520 ;
      RECT 1.7990 0.3490 2.0010 0.3990 ;
      RECT 1.9510 0.3990 2.0010 0.5370 ;
      RECT 1.7990 0.3990 1.8490 1.1020 ;
      RECT 3.9870 1.5280 4.6770 1.5780 ;
      RECT 4.8580 0.6270 5.1330 0.6540 ;
      RECT 4.4430 0.6040 5.1330 0.6270 ;
      RECT 4.4430 0.5770 4.9080 0.6040 ;
      RECT 1.2910 0.3190 1.3930 0.3690 ;
      RECT 1.3430 0.3690 1.3930 1.0020 ;
      RECT 1.2910 0.1510 1.3410 0.3190 ;
      RECT 1.2910 0.1010 1.9410 0.1510 ;
      RECT 0.7190 0.3010 1.1050 0.3510 ;
      RECT 1.4030 0.2040 1.7890 0.2540 ;
      RECT 0.7350 1.3160 1.0890 1.3660 ;
      RECT 0.7350 0.9800 0.7850 1.3160 ;
      RECT 1.0390 1.1920 1.0890 1.3160 ;
      RECT 1.7070 1.4160 1.9460 1.4660 ;
      RECT 2.1630 0.1040 3.0050 0.1540 ;
      RECT 2.7870 0.1540 2.8370 0.2170 ;
      RECT 2.9230 1.4170 3.3090 1.4670 ;
      RECT 2.5590 0.7260 2.6610 0.7760 ;
      RECT 2.5590 0.7760 2.6090 1.1520 ;
      RECT 2.6110 0.6760 2.6610 0.7260 ;
      RECT 2.6110 0.6260 2.7010 0.6760 ;
      RECT 2.6110 0.4960 2.6610 0.6260 ;
      RECT 2.5430 0.4460 2.6610 0.4960 ;
      RECT 5.2030 0.6040 5.4370 0.6540 ;
      RECT 3.9270 0.3000 3.9770 1.2160 ;
      RECT 4.3430 0.5270 4.3930 0.6540 ;
      RECT 4.1390 0.6540 4.3930 0.6770 ;
      RECT 4.1390 0.6770 4.4730 0.7040 ;
      RECT 4.3430 0.7040 4.4730 0.7270 ;
      RECT 4.4230 0.7270 4.4730 1.2160 ;
      RECT 3.9270 1.2160 4.4730 1.2660 ;
      RECT 5.2030 0.5270 5.2530 0.6040 ;
      RECT 4.3430 0.4770 5.2530 0.5270 ;
      RECT 0.7000 0.5730 0.8770 0.6230 ;
      RECT 0.7000 0.6230 0.7500 0.8080 ;
      RECT 0.4310 0.8080 0.7500 0.8580 ;
      RECT 0.4310 0.8580 0.4810 1.2460 ;
      RECT 0.4310 0.4550 0.4810 0.6010 ;
      RECT 0.4710 0.6510 0.5210 0.8080 ;
      RECT 0.4310 0.6010 0.5210 0.6510 ;
  END
END SDFFSSRX2_LVT

MACRO SDFFX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.168 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.9610 1.1610 5.0710 1.2210 ;
        RECT 5.0210 0.2040 5.0710 1.1610 ;
        RECT 4.8390 1.2210 5.0710 1.2710 ;
        RECT 4.8230 0.1540 5.0710 0.2040 ;
        RECT 4.8390 1.2710 4.8890 1.5460 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8090 1.0090 4.9190 1.1190 ;
        RECT 4.8690 0.8540 4.9190 1.0090 ;
        RECT 4.5350 0.8040 4.9190 0.8540 ;
        RECT 4.5350 0.8540 4.5850 1.5460 ;
        RECT 4.8690 0.3590 4.9190 0.8040 ;
        RECT 4.5350 0.3090 4.9190 0.3590 ;
        RECT 4.5350 0.1480 4.5850 0.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7690 1.4240 1.9410 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 5.1680 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 4.6870 1.0190 4.7370 1.6420 ;
        RECT 1.6470 1.1340 1.6970 1.6420 ;
        RECT 4.4230 1.3580 4.4730 1.6420 ;
        RECT 3.8550 1.3580 3.9050 1.6420 ;
        RECT 3.1910 1.3280 3.2410 1.6420 ;
        RECT 2.1030 1.3540 2.1530 1.6420 ;
        RECT 4.3650 1.3080 4.4730 1.3580 ;
        RECT 3.8550 1.3080 3.9930 1.3580 ;
        RECT 2.9980 1.2780 3.2410 1.3280 ;
        RECT 1.9510 1.3040 2.1530 1.3540 ;
        RECT 1.9510 1.0880 2.0010 1.3040 ;
        RECT 2.1030 1.0880 2.1530 1.3040 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 0.6640 1.0110 0.8150 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6800 0.7250 0.7300 ;
        RECT 0.4010 0.5530 0.5110 0.6800 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2360 1.3150 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 5.1680 0.0300 ;
        RECT 1.6470 0.0300 1.6970 0.1960 ;
        RECT 3.0150 0.0300 3.0650 0.1990 ;
        RECT 4.6870 0.0300 4.7370 0.2200 ;
        RECT 0.5830 0.0300 0.6330 0.5150 ;
        RECT 0.4310 0.0300 0.4810 0.4370 ;
        RECT 4.3830 0.0300 4.4330 0.3300 ;
        RECT 1.6470 0.1960 2.1530 0.2460 ;
        RECT 3.0150 0.1990 3.2400 0.2490 ;
        RECT 3.9110 0.3300 4.4490 0.3800 ;
        RECT 2.1030 0.2460 2.1530 0.4500 ;
        RECT 1.9510 0.2460 2.0010 0.4500 ;
        RECT 1.6470 0.2460 1.6970 0.4080 ;
        RECT 3.0150 0.2490 3.0650 0.3730 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 5.2830 1.7730 ;
    LAYER M1 ;
      RECT 3.0910 1.4280 3.1410 1.5840 ;
      RECT 2.4830 1.3780 3.1410 1.4280 ;
      RECT 2.4830 1.4280 2.5330 1.5260 ;
      RECT 2.3150 1.5260 2.5330 1.5760 ;
      RECT 2.6350 1.4780 3.0050 1.5280 ;
      RECT 2.6350 1.5280 2.6850 1.5650 ;
      RECT 3.9860 1.5210 4.3730 1.5710 ;
      RECT 2.9230 0.7580 3.4450 0.8080 ;
      RECT 3.3950 0.5870 3.4450 0.7580 ;
      RECT 2.5590 0.6400 3.3090 0.6900 ;
      RECT 2.5590 0.4840 2.6090 0.6400 ;
      RECT 2.5590 0.6900 2.6090 1.1580 ;
      RECT 2.5590 0.4340 2.7770 0.4840 ;
      RECT 2.5590 1.1580 2.7770 1.2080 ;
      RECT 2.5590 0.3550 2.6090 0.4340 ;
      RECT 2.5590 1.2080 2.6090 1.3140 ;
      RECT 2.4070 0.2990 2.4970 0.3810 ;
      RECT 2.4310 0.3810 2.4810 0.9880 ;
      RECT 2.4070 1.0380 2.4570 1.3140 ;
      RECT 1.0230 0.9880 2.4810 1.0380 ;
      RECT 1.3430 0.4620 1.3930 0.5040 ;
      RECT 1.0230 0.4120 1.3930 0.4620 ;
      RECT 1.6500 0.7760 1.7000 0.9880 ;
      RECT 1.6500 0.7260 1.7370 0.7760 ;
      RECT 1.6870 0.5540 1.7370 0.7260 ;
      RECT 1.3430 0.5040 1.7370 0.5540 ;
      RECT 4.7630 0.4880 4.8130 0.7040 ;
      RECT 3.6230 0.4380 4.8130 0.4880 ;
      RECT 4.4230 0.7040 4.8130 0.7540 ;
      RECT 4.4230 0.7540 4.4730 1.2080 ;
      RECT 4.0630 1.2080 4.4730 1.2580 ;
      RECT 3.6230 0.4880 3.6730 1.1650 ;
      RECT 3.9260 0.4880 3.9760 0.6990 ;
      RECT 3.8350 0.6990 3.9760 0.7490 ;
      RECT 4.0030 0.0880 4.0530 0.2300 ;
      RECT 3.3310 0.2300 4.0530 0.2800 ;
      RECT 3.5310 0.1780 3.6130 0.2300 ;
      RECT 3.3310 0.2800 3.3810 0.3140 ;
      RECT 3.1800 0.3140 3.3810 0.3640 ;
      RECT 3.1800 0.3640 3.2300 0.5400 ;
      RECT 2.9230 0.5400 3.2300 0.5900 ;
      RECT 2.7660 1.0010 3.5610 1.0510 ;
      RECT 3.5110 0.4700 3.5610 1.0010 ;
      RECT 3.4710 1.0510 3.5210 1.3080 ;
      RECT 3.2880 0.4200 3.5610 0.4700 ;
      RECT 3.3190 1.3080 3.5210 1.3580 ;
      RECT 3.4710 0.3710 3.5210 0.4200 ;
      RECT 3.3190 1.1660 3.3690 1.3080 ;
      RECT 1.4520 0.6040 1.6370 0.6540 ;
      RECT 0.2050 0.5280 0.2550 0.8880 ;
      RECT 0.2790 0.9380 0.3290 1.2160 ;
      RECT 0.2050 0.4780 0.3290 0.5280 ;
      RECT 0.2790 0.3180 0.3290 0.4780 ;
      RECT 0.2050 0.8880 1.5020 0.9380 ;
      RECT 1.4520 0.6540 1.5020 0.8880 ;
      RECT 0.8870 0.3120 1.5450 0.3620 ;
      RECT 1.4950 0.3620 1.5450 0.3940 ;
      RECT 0.8870 0.3620 0.9370 0.3940 ;
      RECT 0.7190 0.5120 1.2570 0.5620 ;
      RECT 0.7350 1.0420 0.9370 1.0920 ;
      RECT 0.7350 1.0920 0.7850 1.2160 ;
      RECT 0.8870 1.0920 0.9370 1.2160 ;
      RECT 1.1750 1.0880 1.5610 1.1380 ;
      RECT 2.0110 0.0960 2.7070 0.1460 ;
      RECT 1.7990 0.6180 2.2450 0.6680 ;
      RECT 1.7990 0.6680 1.8490 0.9140 ;
      RECT 1.7990 0.4220 1.8490 0.6180 ;
      RECT 2.2550 0.5180 2.3810 0.5680 ;
      RECT 2.2550 0.3940 2.3050 0.5180 ;
      RECT 2.3310 0.5680 2.3810 0.7180 ;
      RECT 2.2550 0.7180 2.3810 0.7680 ;
      RECT 2.2550 0.7680 2.3050 0.9140 ;
      RECT 4.0400 0.6040 4.6770 0.6540 ;
      RECT 4.0400 0.6540 4.0900 0.9780 ;
      RECT 3.7350 0.9780 4.0900 1.0270 ;
      RECT 3.7350 0.5880 3.7850 0.9780 ;
      RECT 3.7580 1.0270 4.0900 1.0280 ;
      RECT 3.7350 0.5380 3.8650 0.5880 ;
      RECT 4.0400 1.0280 4.0900 1.0290 ;
      RECT 4.1500 0.7090 4.3730 0.7590 ;
      RECT 3.7470 1.1490 3.7970 1.2720 ;
      RECT 3.5710 1.2720 3.7970 1.3220 ;
      RECT 3.5710 1.3220 3.6210 1.5220 ;
      RECT 3.3790 1.5220 3.6210 1.5720 ;
      RECT 4.1500 0.7590 4.2000 1.0990 ;
      RECT 3.7470 1.0990 4.2000 1.1490 ;
    LAYER PO ;
      RECT 3.5570 0.8820 3.5870 1.6060 ;
      RECT 2.9490 0.0680 2.9790 0.6180 ;
      RECT 4.3170 0.0680 4.3470 0.7870 ;
      RECT 2.4930 0.9900 2.5230 1.6060 ;
      RECT 5.0770 0.0680 5.1070 1.6060 ;
      RECT 2.4930 0.0680 2.5230 0.5420 ;
      RECT 4.6210 0.0680 4.6510 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 4.7730 0.0680 4.8030 1.6060 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 3.7090 0.0680 3.7390 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 4.9250 0.0680 4.9550 1.6060 ;
      RECT 4.4690 0.0680 4.4990 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 2.9490 0.7300 2.9790 1.6060 ;
      RECT 3.5570 0.0680 3.5870 0.6220 ;
      RECT 4.3170 1.0120 4.3470 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
  END
END SDFFX1_LVT

MACRO SDFFX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.472 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6870 0.1480 4.7370 0.3940 ;
        RECT 4.6870 0.3940 5.2330 0.4440 ;
        RECT 5.1130 0.4440 5.2330 0.5110 ;
        RECT 5.1830 0.5110 5.2330 0.8040 ;
        RECT 4.6870 0.8040 5.2330 0.8540 ;
        RECT 4.6870 0.8540 4.7370 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7690 1.4240 1.9410 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 5.4720 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 4.8390 0.9600 4.8890 1.6420 ;
        RECT 4.5350 0.8520 4.5850 1.6420 ;
        RECT 1.6470 1.1340 1.6970 1.6420 ;
        RECT 5.1430 1.0520 5.1930 1.6420 ;
        RECT 4.4230 1.3580 4.4730 1.6420 ;
        RECT 3.8550 1.3580 3.9050 1.6420 ;
        RECT 3.1910 1.3280 3.2410 1.6420 ;
        RECT 2.1030 1.3540 2.1530 1.6420 ;
        RECT 4.3650 1.3080 4.4730 1.3580 ;
        RECT 3.8550 1.3080 3.9930 1.3580 ;
        RECT 2.9980 1.2780 3.2410 1.3280 ;
        RECT 1.9510 1.3040 2.1530 1.3540 ;
        RECT 1.9510 1.0880 2.0010 1.3040 ;
        RECT 2.1030 1.0880 2.1530 1.3040 ;
    END
  END VDD

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2650 0.0970 5.3750 0.2070 ;
        RECT 5.3070 0.2070 5.3570 0.2700 ;
        RECT 4.9910 0.2700 5.3570 0.3200 ;
        RECT 4.9910 0.1480 5.0410 0.2700 ;
        RECT 5.3070 0.3200 5.3570 0.9180 ;
        RECT 4.9910 0.9180 5.3570 0.9680 ;
        RECT 4.9910 0.9680 5.0410 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 0.6640 1.0110 0.8150 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6800 0.7250 0.7300 ;
        RECT 0.4010 0.5530 0.5110 0.6800 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2360 1.3150 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 5.4720 0.0300 ;
        RECT 1.6470 0.0300 1.6970 0.1960 ;
        RECT 3.0150 0.0300 3.0650 0.1990 ;
        RECT 0.5830 0.0300 0.6330 0.5150 ;
        RECT 0.4310 0.0300 0.4810 0.4370 ;
        RECT 5.1430 0.0300 5.1930 0.2200 ;
        RECT 4.8390 0.0300 4.8890 0.3190 ;
        RECT 4.5350 0.0300 4.5850 0.4080 ;
        RECT 4.3830 0.0300 4.4330 0.3300 ;
        RECT 1.6470 0.1960 2.1530 0.2460 ;
        RECT 3.0150 0.1990 3.2400 0.2490 ;
        RECT 3.9110 0.3300 4.4490 0.3800 ;
        RECT 2.1030 0.2460 2.1530 0.4500 ;
        RECT 1.9510 0.2460 2.0010 0.4500 ;
        RECT 1.6470 0.2460 1.6970 0.4080 ;
        RECT 3.0150 0.2490 3.0650 0.3730 ;
    END
  END VSS
  OBS
    LAYER PO ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 2.9490 0.7300 2.9790 1.6060 ;
      RECT 3.5570 0.0680 3.5870 0.6220 ;
      RECT 4.3170 1.0120 4.3470 1.6060 ;
      RECT 5.3810 0.0680 5.4110 1.6060 ;
      RECT 5.0770 0.0680 5.1070 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 5.2290 0.0680 5.2590 1.6060 ;
      RECT 3.5570 0.8820 3.5870 1.6060 ;
      RECT 2.9490 0.0680 2.9790 0.6180 ;
      RECT 4.3170 0.0680 4.3470 0.7870 ;
      RECT 2.4930 0.9900 2.5230 1.6060 ;
      RECT 2.4930 0.0680 2.5230 0.5420 ;
      RECT 4.6210 0.0680 4.6510 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 4.7730 0.0680 4.8030 1.6060 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 3.7090 0.0680 3.7390 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 4.9250 0.0680 4.9550 1.6060 ;
      RECT 4.4690 0.0680 4.4990 1.6060 ;
    LAYER NWELL ;
      RECT -0.1150 0.6790 5.5870 1.7730 ;
    LAYER M1 ;
      RECT 4.0030 0.0880 4.0530 0.2300 ;
      RECT 3.3310 0.2300 4.0530 0.2800 ;
      RECT 3.5310 0.1780 3.6130 0.2300 ;
      RECT 3.3310 0.2800 3.3810 0.3140 ;
      RECT 3.1800 0.3140 3.3810 0.3640 ;
      RECT 3.1800 0.3640 3.2300 0.5400 ;
      RECT 2.9230 0.5400 3.2300 0.5900 ;
      RECT 2.7660 1.0010 3.5610 1.0510 ;
      RECT 3.5110 0.4700 3.5610 1.0010 ;
      RECT 3.4710 1.0510 3.5210 1.3080 ;
      RECT 3.2880 0.4200 3.5610 0.4700 ;
      RECT 3.3190 1.3080 3.5210 1.3580 ;
      RECT 3.4710 0.3710 3.5210 0.4200 ;
      RECT 3.3190 1.1660 3.3690 1.3080 ;
      RECT 1.4520 0.6040 1.6370 0.6540 ;
      RECT 0.2050 0.5280 0.2550 0.8880 ;
      RECT 0.2790 0.9380 0.3290 1.2160 ;
      RECT 0.2050 0.4780 0.3290 0.5280 ;
      RECT 0.2790 0.3180 0.3290 0.4780 ;
      RECT 0.2050 0.8880 1.5020 0.9380 ;
      RECT 1.4520 0.6540 1.5020 0.8880 ;
      RECT 0.7350 1.0420 0.9370 1.0920 ;
      RECT 0.7350 1.0920 0.7850 1.2160 ;
      RECT 0.8870 1.0920 0.9370 1.2160 ;
      RECT 1.1750 1.0880 1.5610 1.1380 ;
      RECT 0.8870 0.3120 1.5450 0.3620 ;
      RECT 0.8870 0.3620 0.9370 0.3940 ;
      RECT 1.4950 0.3620 1.5450 0.3940 ;
      RECT 2.0110 0.0960 2.7070 0.1460 ;
      RECT 1.7990 0.6180 2.2450 0.6680 ;
      RECT 1.7990 0.6680 1.8490 0.9140 ;
      RECT 1.7990 0.4220 1.8490 0.6180 ;
      RECT 2.2550 0.5180 2.3810 0.5680 ;
      RECT 2.2550 0.3940 2.3050 0.5180 ;
      RECT 2.3310 0.5680 2.3810 0.7180 ;
      RECT 2.2550 0.7180 2.3810 0.7680 ;
      RECT 2.2550 0.7680 2.3050 0.9140 ;
      RECT 4.0400 0.6040 4.8290 0.6540 ;
      RECT 4.0400 0.6540 4.0900 0.9780 ;
      RECT 3.7350 0.9780 4.0900 1.0270 ;
      RECT 3.7350 0.5880 3.7850 0.9780 ;
      RECT 3.7580 1.0270 4.0900 1.0280 ;
      RECT 3.7350 0.5380 3.8650 0.5880 ;
      RECT 4.0400 1.0280 4.0900 1.0290 ;
      RECT 4.1500 0.7090 4.3730 0.7590 ;
      RECT 3.7470 1.1490 3.7970 1.2720 ;
      RECT 3.5710 1.2720 3.7970 1.3220 ;
      RECT 3.5710 1.3220 3.6210 1.5220 ;
      RECT 3.3790 1.5220 3.6210 1.5720 ;
      RECT 4.1500 0.7590 4.2000 1.0990 ;
      RECT 3.7470 1.0990 4.2000 1.1490 ;
      RECT 2.3150 1.5260 2.5330 1.5760 ;
      RECT 2.4830 1.4280 2.5330 1.5260 ;
      RECT 2.4830 1.3780 3.1410 1.4280 ;
      RECT 3.0910 1.4280 3.1410 1.5840 ;
      RECT 2.6350 1.4780 3.0050 1.5280 ;
      RECT 2.6350 1.5280 2.6850 1.5650 ;
      RECT 3.9860 1.5210 4.3730 1.5710 ;
      RECT 0.7190 0.5120 1.2570 0.5620 ;
      RECT 2.9230 0.7580 3.4450 0.8080 ;
      RECT 3.3950 0.5870 3.4450 0.7580 ;
      RECT 2.5590 0.6400 3.3090 0.6900 ;
      RECT 2.5590 0.4840 2.6090 0.6400 ;
      RECT 2.5590 0.6900 2.6090 1.1580 ;
      RECT 2.5590 0.4340 2.7770 0.4840 ;
      RECT 2.5590 1.1580 2.7770 1.2080 ;
      RECT 2.5590 0.3550 2.6090 0.4340 ;
      RECT 2.5590 1.2080 2.6090 1.3140 ;
      RECT 2.4070 0.2990 2.4970 0.3810 ;
      RECT 2.4310 0.3810 2.4810 0.9880 ;
      RECT 2.4070 1.0380 2.4570 1.3140 ;
      RECT 1.0230 0.9880 2.4810 1.0380 ;
      RECT 1.3430 0.4620 1.3930 0.5040 ;
      RECT 1.0230 0.4120 1.3930 0.4620 ;
      RECT 1.6500 0.7760 1.7000 0.9880 ;
      RECT 1.6500 0.7260 1.7370 0.7760 ;
      RECT 1.6870 0.5540 1.7370 0.7260 ;
      RECT 1.3430 0.5040 1.7370 0.5540 ;
      RECT 4.8960 0.6040 5.1330 0.6540 ;
      RECT 4.8960 0.6540 4.9460 0.7040 ;
      RECT 4.8960 0.5440 4.9460 0.6040 ;
      RECT 4.4330 0.7040 4.9460 0.7540 ;
      RECT 3.9260 0.4940 4.9460 0.5440 ;
      RECT 4.4340 0.7540 4.4840 1.2080 ;
      RECT 3.9260 0.5440 3.9760 0.6990 ;
      RECT 3.9260 0.4880 3.9760 0.4940 ;
      RECT 4.0630 1.2080 4.4840 1.2580 ;
      RECT 3.8350 0.6990 3.9760 0.7490 ;
      RECT 3.6230 0.4380 3.9760 0.4880 ;
      RECT 3.6230 0.4880 3.6730 1.1650 ;
  END
END SDFFX2_LVT

MACRO SHFILL128_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 19.456 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 19.4560 1.7020 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 19.4560 0.0300 ;
    END
  END VSS
  OBS
    LAYER PO ;
      RECT 3.7090 0.0660 3.7390 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 9.7890 0.0660 9.8190 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 19.3650 0.0660 19.3950 1.6060 ;
      RECT 18.7570 0.0660 18.7870 1.6060 ;
      RECT 18.6050 0.0660 18.6350 1.6060 ;
      RECT 18.4530 0.0660 18.4830 1.6060 ;
      RECT 18.3010 0.0660 18.3310 1.6060 ;
      RECT 16.3250 0.0660 16.3550 1.6060 ;
      RECT 16.1730 0.0660 16.2030 1.6060 ;
      RECT 16.0210 0.0660 16.0510 1.6060 ;
      RECT 15.8690 0.0660 15.8990 1.6060 ;
      RECT 13.5890 0.0660 13.6190 1.6060 ;
      RECT 13.4370 0.0660 13.4670 1.6060 ;
      RECT 13.7410 0.0660 13.7710 1.6060 ;
      RECT 13.8930 0.0660 13.9230 1.6060 ;
      RECT 14.5010 0.0660 14.5310 1.6060 ;
      RECT 14.3490 0.0660 14.3790 1.6060 ;
      RECT 14.1970 0.0660 14.2270 1.6060 ;
      RECT 14.0450 0.0660 14.0750 1.6060 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 10.8530 0.0660 10.8830 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 11.3090 0.0660 11.3390 1.6060 ;
      RECT 11.4610 0.0660 11.4910 1.6060 ;
      RECT 13.1330 0.0660 13.1630 1.6060 ;
      RECT 13.2850 0.0660 13.3150 1.6060 ;
      RECT 12.6770 0.0660 12.7070 1.6060 ;
      RECT 12.5250 0.0660 12.5550 1.6060 ;
      RECT 12.3730 0.0660 12.4030 1.6060 ;
      RECT 10.2450 0.0660 10.2750 1.6060 ;
      RECT 10.0930 0.0660 10.1230 1.6060 ;
      RECT 9.9410 0.0660 9.9710 1.6060 ;
      RECT 16.9330 0.0660 16.9630 1.6060 ;
      RECT 16.7810 0.0660 16.8110 1.6060 ;
      RECT 16.6290 0.0660 16.6590 1.6060 ;
      RECT 16.4770 0.0660 16.5070 1.6060 ;
      RECT 15.2610 0.0660 15.2910 1.6060 ;
      RECT 15.4130 0.0660 15.4430 1.6060 ;
      RECT 15.5650 0.0660 15.5950 1.6060 ;
      RECT 15.7170 0.0660 15.7470 1.6060 ;
      RECT 15.1090 0.0660 15.1390 1.6060 ;
      RECT 14.9570 0.0660 14.9870 1.6060 ;
      RECT 14.8050 0.0660 14.8350 1.6060 ;
      RECT 14.6530 0.0660 14.6830 1.6060 ;
      RECT 11.9170 0.0660 11.9470 1.6060 ;
      RECT 12.0690 0.0660 12.0990 1.6060 ;
      RECT 17.0850 0.0660 17.1150 1.6060 ;
      RECT 12.2210 0.0660 12.2510 1.6060 ;
      RECT 17.2370 0.0660 17.2670 1.6060 ;
      RECT 17.3890 0.0660 17.4190 1.6060 ;
      RECT 17.5410 0.0660 17.5710 1.6060 ;
      RECT 18.1490 0.0660 18.1790 1.6060 ;
      RECT 17.9970 0.0660 18.0270 1.6060 ;
      RECT 17.8450 0.0660 17.8750 1.6060 ;
      RECT 17.6930 0.0660 17.7230 1.6060 ;
      RECT 18.9090 0.0660 18.9390 1.6060 ;
      RECT 19.0610 0.0660 19.0910 1.6060 ;
      RECT 19.2130 0.0660 19.2430 1.6060 ;
      RECT 11.1570 0.0660 11.1870 1.6060 ;
      RECT 11.0050 0.0660 11.0350 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 9.3330 0.0660 9.3630 1.6060 ;
      RECT 9.4850 0.0660 9.5150 1.6060 ;
      RECT 9.6370 0.0660 9.6670 1.6060 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 12.9810 0.0660 13.0110 1.6060 ;
      RECT 12.8290 0.0660 12.8590 1.6060 ;
      RECT 11.7650 0.0660 11.7950 1.6060 ;
      RECT 11.6130 0.0660 11.6430 1.6060 ;
      RECT 10.3970 0.0660 10.4270 1.6060 ;
      RECT 10.5490 0.0660 10.5790 1.6060 ;
      RECT 10.7010 0.0660 10.7310 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
    LAYER NWELL ;
      RECT -0.1150 0.6790 19.5710 1.7730 ;
  END
END SHFILL128_LVT

MACRO SHFILL1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.152 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 0.1520 1.7020 ;
        RECT 0.0510 1.6240 0.1010 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 0.1520 0.0300 ;
        RECT 0.0510 0.0300 0.1010 0.0480 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1490 0.6790 0.3010 1.7730 ;
    LAYER PO ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
  END
END SHFILL1_LVT

MACRO SHFILL2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.304 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 0.3040 1.7020 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 0.3040 0.0300 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 0.4190 1.7730 ;
    LAYER PO ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
  END
END SHFILL2_LVT

MACRO SHFILL3_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.456 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 0.4560 1.7020 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 0.4560 0.0300 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 0.5710 1.7730 ;
    LAYER PO ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
  END
END SHFILL3_LVT

MACRO SHFILL64_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.728 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 9.7280 1.7020 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 9.7280 0.0300 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 9.8430 1.7730 ;
    LAYER PO ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 9.3330 0.0660 9.3630 1.6060 ;
      RECT 9.4850 0.0660 9.5150 1.6060 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 9.6370 0.0660 9.6670 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 3.7090 0.0660 3.7390 1.6060 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
  END
END SHFILL64_LVT

MACRO TIEH_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.76 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 1.1610 0.5140 1.2740 ;
        RECT 0.4310 1.2740 0.4810 1.5490 ;
        RECT 0.4310 0.8230 0.4810 1.1610 ;
    END
    ANTENNADIFFAREA 0.0816 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.2490 1.3130 0.3620 1.4230 ;
        RECT 0.2790 0.8230 0.3290 1.3130 ;
        RECT 0.2790 1.4230 0.3290 1.6420 ;
        RECT 0.0000 1.6420 0.7600 1.7020 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 0.7600 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.5390 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 0.8750 1.7730 ;
    LAYER M1 ;
      RECT 0.4310 0.1910 0.4810 0.6970 ;
      RECT 0.3390 0.6470 0.4810 0.6970 ;
    LAYER PO ;
      RECT 0.3650 0.0690 0.3950 1.6060 ;
      RECT 0.2130 0.0710 0.2430 1.6060 ;
      RECT 0.6690 0.0710 0.6990 1.6060 ;
      RECT 0.5170 0.0710 0.5470 1.6060 ;
      RECT 0.0610 0.0710 0.0910 1.6060 ;
  END
END TIEH_LVT

MACRO TIEL_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.76 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 0.2490 0.5140 0.3590 ;
        RECT 0.4310 0.3590 0.4810 0.6100 ;
        RECT 0.4310 0.2450 0.4810 0.2490 ;
    END
    ANTENNADIFFAREA 0.0428 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 0.7600 1.7020 ;
        RECT 0.2790 0.8230 0.3290 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 0.7600 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.4010 ;
        RECT 0.2490 0.4010 0.3620 0.5110 ;
        RECT 0.2790 0.5110 0.3290 0.5390 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 0.8750 1.7730 ;
    LAYER M1 ;
      RECT 0.4310 0.6850 0.4810 1.5490 ;
      RECT 0.3390 0.6600 0.4810 0.7100 ;
    LAYER PO ;
      RECT 0.3650 0.0690 0.3950 1.6060 ;
      RECT 0.2130 0.0710 0.2430 1.6060 ;
      RECT 0.6690 0.0710 0.6990 1.6060 ;
      RECT 0.5170 0.0710 0.5470 1.6060 ;
      RECT 0.0610 0.0710 0.0910 1.6060 ;
  END
END TIEL_LVT

MACRO TNBUFFX16_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.168 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4360 1.3710 1.0400 1.4210 ;
        RECT 0.5530 1.4210 0.6630 1.4230 ;
        RECT 0.5530 1.3130 0.6630 1.3710 ;
        RECT 0.4360 1.1440 0.4860 1.3710 ;
        RECT 0.3310 1.0940 0.4860 1.1440 ;
        RECT 0.3310 0.7100 0.3810 1.0940 ;
        RECT 0.3310 0.6600 0.4210 0.7100 ;
    END
    ANTENNAGATEAREA 0.0753 ;
  END EN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 5.1680 1.7020 ;
        RECT 4.6870 1.2720 4.7370 1.6420 ;
        RECT 4.3830 1.2720 4.4330 1.6420 ;
        RECT 4.0790 1.2720 4.1290 1.6420 ;
        RECT 3.7750 1.2720 3.8250 1.6420 ;
        RECT 3.4710 1.2720 3.5210 1.6420 ;
        RECT 3.1670 1.2720 3.2170 1.6420 ;
        RECT 2.8630 1.2720 2.9130 1.6420 ;
        RECT 0.2790 1.2140 0.3290 1.6420 ;
        RECT 2.5590 1.2750 2.6090 1.6420 ;
        RECT 1.1910 1.3210 1.2410 1.6420 ;
        RECT 0.7350 1.2710 1.5450 1.3210 ;
        RECT 0.7350 1.0900 0.7850 1.2710 ;
        RECT 1.1910 1.0900 1.2410 1.2710 ;
        RECT 1.0390 1.0900 1.0890 1.2710 ;
        RECT 1.4950 1.0900 1.5450 1.2710 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 5.1680 0.0300 ;
        RECT 2.8630 0.0300 2.9130 0.3680 ;
        RECT 4.6870 0.0300 4.7370 0.3680 ;
        RECT 4.3830 0.0300 4.4330 0.3680 ;
        RECT 4.0790 0.0300 4.1290 0.3680 ;
        RECT 3.7750 0.0300 3.8250 0.3680 ;
        RECT 3.4710 0.0300 3.5210 0.3680 ;
        RECT 3.1670 0.0300 3.2170 0.3680 ;
        RECT 0.2790 0.0300 0.3290 0.5740 ;
        RECT 2.5590 0.0300 2.6090 0.2150 ;
        RECT 1.3430 0.2150 2.6090 0.2650 ;
        RECT 1.8000 0.2650 1.8500 0.4320 ;
        RECT 1.3430 0.2650 1.3930 0.4450 ;
        RECT 1.6470 0.2650 1.6970 0.4330 ;
        RECT 2.1040 0.2650 2.1540 0.4330 ;
        RECT 2.5590 0.2650 2.6090 0.3680 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.9270 1.1340 3.9770 1.4720 ;
        RECT 4.2310 1.1340 4.2810 1.4720 ;
        RECT 4.5350 1.1340 4.5850 1.4720 ;
        RECT 4.8390 1.1340 4.8890 1.4720 ;
        RECT 2.4070 1.1340 2.4570 1.4720 ;
        RECT 2.7110 1.1340 2.7610 1.4720 ;
        RECT 3.0150 1.1340 3.0650 1.4720 ;
        RECT 3.3190 1.1340 3.3690 1.4720 ;
        RECT 3.6230 1.1340 3.6730 1.4720 ;
        RECT 2.4070 1.0840 4.9610 1.1340 ;
        RECT 3.9270 0.9000 3.9770 1.0840 ;
        RECT 4.2310 0.9000 4.2810 1.0840 ;
        RECT 4.5350 0.9000 4.5850 1.0840 ;
        RECT 2.7110 0.9000 2.7610 1.0840 ;
        RECT 3.0150 0.9000 3.0650 1.0840 ;
        RECT 3.3190 0.9000 3.3690 1.0840 ;
        RECT 3.6230 0.9000 3.6730 1.0840 ;
        RECT 4.9110 0.6630 4.9610 1.0840 ;
        RECT 4.9110 0.5530 5.0710 0.6630 ;
        RECT 4.9110 0.4890 4.9610 0.5530 ;
        RECT 4.8390 0.4880 4.9610 0.4890 ;
        RECT 2.4070 0.4390 4.9610 0.4880 ;
        RECT 2.4070 0.4380 4.9130 0.4390 ;
        RECT 2.7110 0.1420 2.7610 0.4380 ;
        RECT 3.0150 0.1420 3.0650 0.4380 ;
        RECT 3.3190 0.1420 3.3690 0.4380 ;
        RECT 3.6230 0.1420 3.6730 0.4380 ;
        RECT 2.4070 0.3910 2.4570 0.4380 ;
        RECT 3.9270 0.1420 3.9770 0.4380 ;
        RECT 4.2310 0.1420 4.2810 0.4380 ;
        RECT 4.5350 0.1420 4.5850 0.4380 ;
        RECT 4.8390 0.1550 4.8890 0.4380 ;
    END
    ANTENNADIFFAREA 1.1532 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 0.6510 1.6520 0.7010 ;
        RECT 1.1610 0.7010 1.2710 0.8150 ;
    END
    ANTENNAGATEAREA 0.1098 ;
  END A
  OBS
    LAYER NWELL ;
      RECT -0.1120 0.6790 5.2800 1.7730 ;
    LAYER M1 ;
      RECT 2.4520 0.7450 4.8440 0.7950 ;
      RECT 1.3430 1.0340 1.3930 1.2020 ;
      RECT 1.3430 0.8000 1.3930 0.9840 ;
      RECT 1.6470 1.0340 1.6970 1.4780 ;
      RECT 1.6470 0.8000 1.6970 0.9840 ;
      RECT 1.8000 1.0340 1.8500 1.2020 ;
      RECT 2.1040 1.0340 2.1540 1.2020 ;
      RECT 2.4830 0.7950 2.5330 0.9840 ;
      RECT 0.5830 0.9840 2.5330 1.0340 ;
      RECT 0.5830 1.0340 0.6330 1.2110 ;
      RECT 0.5830 0.2830 0.6330 0.9840 ;
      RECT 0.8870 1.0340 0.9370 1.2110 ;
      RECT 0.8870 0.3090 0.9370 0.9840 ;
      RECT 0.4310 0.1000 2.2600 0.1500 ;
      RECT 0.4310 0.1500 0.4810 0.5600 ;
      RECT 0.4310 0.7890 0.5210 0.8400 ;
      RECT 0.4310 0.8400 0.4810 1.0160 ;
      RECT 0.4310 0.5600 0.5210 0.6100 ;
      RECT 0.4710 0.6100 0.5210 0.7890 ;
      RECT 1.0390 0.5390 4.8440 0.5890 ;
      RECT 1.1910 0.2360 1.2410 0.5390 ;
      RECT 1.4950 0.3280 1.5450 0.5390 ;
      RECT 1.9510 0.3690 2.0010 0.5390 ;
      RECT 1.9510 0.7720 2.0010 0.9110 ;
      RECT 2.2550 0.5890 2.3050 0.7220 ;
      RECT 2.2550 0.3480 2.3050 0.5390 ;
      RECT 1.9510 0.7220 2.3050 0.7720 ;
      RECT 2.2550 0.7720 2.3050 0.9260 ;
      RECT 1.0390 0.2590 1.0890 0.5390 ;
      RECT 0.7350 0.2090 1.0890 0.2590 ;
      RECT 0.7350 0.2590 0.7850 0.5790 ;
    LAYER PO ;
      RECT 3.4050 0.0660 3.4350 0.6170 ;
      RECT 3.4050 0.7170 3.4350 1.6060 ;
      RECT 3.1010 0.0660 3.1310 0.6170 ;
      RECT 3.1010 0.7170 3.1310 1.6060 ;
      RECT 2.6450 0.7170 2.6750 1.6060 ;
      RECT 2.7970 0.7170 2.8270 1.6060 ;
      RECT 2.9490 0.7170 2.9790 1.6060 ;
      RECT 2.4930 0.7170 2.5230 1.6060 ;
      RECT 2.4930 0.0660 2.5230 0.6170 ;
      RECT 2.9490 0.0660 2.9790 0.6170 ;
      RECT 2.7970 0.0660 2.8270 0.6170 ;
      RECT 2.6450 0.0660 2.6750 0.6170 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 4.7730 0.0660 4.8030 0.6170 ;
      RECT 4.7730 0.7170 4.8030 1.6060 ;
      RECT 4.4690 0.0660 4.4990 0.6170 ;
      RECT 4.4690 0.7170 4.4990 1.6060 ;
      RECT 4.3170 0.0660 4.3470 0.6170 ;
      RECT 4.3170 0.7170 4.3470 1.6060 ;
      RECT 4.6210 0.0660 4.6510 0.6170 ;
      RECT 4.6210 0.7170 4.6510 1.6060 ;
      RECT 4.1650 0.0660 4.1950 0.6170 ;
      RECT 4.1650 0.7170 4.1950 1.6060 ;
      RECT 4.0130 0.0660 4.0430 0.6170 ;
      RECT 4.0130 0.7170 4.0430 1.6060 ;
      RECT 3.8610 0.0660 3.8910 0.6170 ;
      RECT 3.8610 0.7170 3.8910 1.6060 ;
      RECT 3.7090 0.0660 3.7390 0.6170 ;
      RECT 3.7090 0.7170 3.7390 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 3.2530 0.0660 3.2830 0.6170 ;
      RECT 3.2530 0.7170 3.2830 1.6060 ;
      RECT 3.5570 0.0660 3.5870 0.6170 ;
      RECT 3.5570 0.7170 3.5870 1.6060 ;
  END
END TNBUFFX16_LVT

MACRO TNBUFFX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.976 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3240 1.3730 0.7360 1.4230 ;
        RECT 0.5530 1.4230 0.6630 1.5750 ;
    END
    ANTENNAGATEAREA 0.0252 ;
  END EN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.9760 1.7020 ;
        RECT 1.4950 1.0840 1.5450 1.6420 ;
        RECT 0.2240 1.2060 0.2740 1.6420 ;
        RECT 0.8100 1.1100 0.8600 1.6420 ;
        RECT 0.2240 1.1560 0.3290 1.2060 ;
        RECT 0.7350 1.0600 0.9370 1.1100 ;
        RECT 0.2790 0.7310 0.3290 1.1560 ;
        RECT 0.7350 0.8140 0.7850 1.0600 ;
        RECT 0.8870 0.8140 0.9370 1.0600 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.9760 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.5420 ;
        RECT 1.4950 0.0300 1.5450 0.2480 ;
        RECT 1.0390 0.2480 1.5450 0.2980 ;
        RECT 1.0390 0.2980 1.0890 0.5520 ;
        RECT 1.1920 0.2980 1.2420 0.5520 ;
        RECT 1.4950 0.2980 1.5450 0.4870 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7020 0.4170 1.7520 0.6780 ;
        RECT 1.7020 0.6780 1.8990 0.8150 ;
        RECT 1.6470 0.3670 1.7520 0.4170 ;
        RECT 1.7020 0.8150 1.7520 1.0840 ;
        RECT 1.6470 0.1030 1.6970 0.3670 ;
        RECT 1.6470 1.0840 1.7520 1.1340 ;
        RECT 1.6470 1.1340 1.6970 1.4720 ;
    END
    ANTENNADIFFAREA 0.1111 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9320 1.4030 1.1190 1.4530 ;
        RECT 1.0090 1.3130 1.1190 1.4030 ;
    END
    ANTENNAGATEAREA 0.0186 ;
  END A
  OBS
    LAYER NWELL ;
      RECT -0.1120 0.6790 2.0880 1.7730 ;
    LAYER M1 ;
      RECT 1.4430 0.5370 1.6520 0.5870 ;
      RECT 1.4430 0.5870 1.4930 0.6020 ;
      RECT 0.8120 0.6020 1.4930 0.6520 ;
      RECT 0.8120 0.5520 0.8620 0.6020 ;
      RECT 0.7350 0.5020 0.9370 0.5520 ;
      RECT 0.8870 0.3480 0.9370 0.5020 ;
      RECT 0.7350 0.3480 0.7850 0.5020 ;
      RECT 1.3430 0.6520 1.3930 0.9340 ;
      RECT 1.3430 0.3480 1.3930 0.6020 ;
      RECT 1.4860 0.7450 1.6520 0.7950 ;
      RECT 1.4860 0.7950 1.5360 0.9840 ;
      RECT 1.4860 0.7440 1.5360 0.7450 ;
      RECT 1.1920 0.9840 1.5360 1.0340 ;
      RECT 0.5830 0.3480 0.6330 0.7140 ;
      RECT 0.5830 0.7640 0.6330 1.0180 ;
      RECT 1.0390 0.7640 1.0890 1.1100 ;
      RECT 1.1920 0.7640 1.2420 0.9840 ;
      RECT 1.1920 0.7130 1.2420 0.7140 ;
      RECT 0.5830 0.7140 1.2420 0.7640 ;
      RECT 0.4310 0.0910 1.3480 0.1410 ;
      RECT 0.4310 0.1410 0.4810 1.1190 ;
    LAYER PO ;
      RECT 1.5810 0.7170 1.6110 1.6060 ;
      RECT 1.5810 0.0640 1.6110 0.6150 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
  END
END TNBUFFX1_LVT

MACRO SDFFASRSX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.232 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2640 0.2340 6.1930 0.2840 ;
        RECT 5.2640 0.2840 5.3750 0.3590 ;
        RECT 6.1430 0.2840 6.1930 1.1560 ;
        RECT 5.7510 1.1560 6.1930 1.2060 ;
        RECT 5.7510 1.2060 5.8010 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4470 1.0500 6.0930 1.1000 ;
        RECT 5.5690 1.1000 5.6870 1.1190 ;
        RECT 5.5690 1.0090 5.6870 1.0500 ;
        RECT 5.4470 1.1000 5.4970 1.5460 ;
        RECT 6.0430 0.3840 6.0930 1.0500 ;
        RECT 5.4280 0.3340 6.0930 0.3840 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 6.2320 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 1.6470 1.1340 1.6970 1.6420 ;
        RECT 5.9030 1.2700 5.9530 1.6420 ;
        RECT 5.2950 1.3630 5.3450 1.6420 ;
        RECT 5.5990 1.2230 5.6490 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 5.0310 1.3580 5.0810 1.6420 ;
        RECT 3.3430 1.3280 3.3930 1.6420 ;
        RECT 2.1030 1.3540 2.1530 1.6420 ;
        RECT 4.2020 1.3080 5.0810 1.3580 ;
        RECT 3.1500 1.2780 3.5520 1.3280 ;
        RECT 1.9510 1.3040 2.1530 1.3540 ;
        RECT 1.9510 1.0880 2.0010 1.3040 ;
        RECT 2.1030 1.1010 2.1530 1.3040 ;
    END
  END VDD

  PIN SO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2650 1.1610 5.3830 1.2710 ;
        RECT 5.2950 0.9270 5.3450 1.1610 ;
        RECT 5.1430 0.8770 5.9930 0.9270 ;
        RECT 5.1430 0.9270 5.1930 1.5460 ;
        RECT 5.9430 0.4840 5.9930 0.8770 ;
        RECT 5.1430 0.4340 5.9930 0.4840 ;
        RECT 5.1430 0.1480 5.1930 0.4340 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END SO

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 0.6640 1.0110 0.8150 ;
    END
    ANTENNAGATEAREA 0.0291 ;
  END D

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.1390 0.1380 4.2210 0.1740 ;
        RECT 2.9390 0.0880 4.2210 0.1380 ;
        RECT 2.9390 0.1380 3.0950 0.2070 ;
    END
    ANTENNAGATEAREA 0.039 ;
  END RSTB

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6800 0.7250 0.7300 ;
        RECT 0.4010 0.5530 0.5110 0.6800 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2360 1.3150 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.7470 0.8460 4.9190 1.0230 ;
    END
    ANTENNAGATEAREA 0.0435 ;
  END SETB

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 6.2320 0.0300 ;
        RECT 1.6470 0.0300 1.6970 0.1960 ;
        RECT 0.5830 0.0300 0.6330 0.5150 ;
        RECT 0.4310 0.0300 0.4810 0.4370 ;
        RECT 2.7570 0.0300 2.8070 0.2870 ;
        RECT 4.9910 0.0300 5.0410 0.3300 ;
        RECT 5.9360 0.0300 5.9860 0.1340 ;
        RECT 1.6470 0.1960 2.1530 0.2460 ;
        RECT 2.7570 0.2870 3.3690 0.3370 ;
        RECT 4.3670 0.3300 5.0570 0.3800 ;
        RECT 5.2760 0.1340 5.9860 0.1840 ;
        RECT 2.1030 0.2460 2.1530 0.4500 ;
        RECT 1.9510 0.2460 2.0010 0.4500 ;
        RECT 1.6470 0.2460 1.6970 0.4080 ;
        RECT 3.3190 0.3370 3.3690 0.4610 ;
        RECT 3.1670 0.3370 3.2170 0.4610 ;
    END
  END VSS

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7690 1.4240 1.9410 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  OBS
    LAYER PO ;
      RECT 2.4930 0.9900 2.5230 1.6060 ;
      RECT 4.9250 0.0680 4.9550 0.7900 ;
      RECT 3.1010 0.0680 3.1310 0.7040 ;
      RECT 3.8610 0.8820 3.8910 1.6060 ;
      RECT 5.3810 0.0680 5.4110 1.6060 ;
      RECT 5.2290 0.0680 5.2590 1.6060 ;
      RECT 5.9890 0.0680 6.0190 1.6060 ;
      RECT 5.8370 0.0680 5.8670 1.6060 ;
      RECT 5.6850 0.0680 5.7150 1.6060 ;
      RECT 5.5330 0.0680 5.5630 1.6060 ;
      RECT 6.1410 0.0680 6.1710 1.6060 ;
      RECT 4.9250 0.9120 4.9550 1.6060 ;
      RECT 3.8610 0.0680 3.8910 0.6220 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 3.1010 0.8260 3.1310 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 4.3170 0.0680 4.3470 1.6060 ;
      RECT 4.7730 0.0680 4.8030 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 3.7090 0.0680 3.7390 1.6060 ;
      RECT 4.4690 0.0680 4.4990 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 4.6210 0.0680 4.6510 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 5.0770 0.0680 5.1070 1.6060 ;
      RECT 2.4930 0.0680 2.5230 0.5420 ;
    LAYER NWELL ;
      RECT -0.1150 0.6790 6.3470 1.7730 ;
    LAYER M1 ;
      RECT 2.4070 1.0380 2.4570 1.3140 ;
      RECT 2.4310 0.3810 2.4810 0.9880 ;
      RECT 2.4070 0.2990 2.4970 0.3810 ;
      RECT 1.0230 0.9880 2.4810 1.0380 ;
      RECT 1.3430 0.4620 1.3930 0.5040 ;
      RECT 1.0230 0.4120 1.3930 0.4620 ;
      RECT 1.6500 0.7760 1.7000 0.9880 ;
      RECT 1.6500 0.7260 1.7370 0.7760 ;
      RECT 1.6870 0.5540 1.7370 0.7260 ;
      RECT 1.3430 0.5040 1.7370 0.5540 ;
      RECT 3.0750 0.8560 3.7650 0.9060 ;
      RECT 5.6560 0.6600 5.8930 0.7100 ;
      RECT 5.6560 0.5840 5.7060 0.6600 ;
      RECT 5.6560 0.7100 5.7060 0.7610 ;
      RECT 4.6780 0.5600 5.7060 0.5840 ;
      RECT 5.0310 0.7610 5.7060 0.8110 ;
      RECT 4.6780 0.5340 5.7020 0.5600 ;
      RECT 5.0310 0.8110 5.0810 1.1080 ;
      RECT 4.6780 0.4880 4.7280 0.5340 ;
      RECT 4.6710 1.1080 5.0810 1.1580 ;
      RECT 4.2300 0.4380 4.7280 0.4880 ;
      RECT 4.2300 0.7660 4.3730 0.8160 ;
      RECT 4.2300 0.4880 4.2800 0.7660 ;
      RECT 4.2300 0.3960 4.2800 0.4380 ;
      RECT 3.9270 0.3460 4.2800 0.3960 ;
      RECT 3.9270 0.3960 3.9770 1.1650 ;
      RECT 3.5020 1.5280 4.8420 1.5780 ;
      RECT 2.3150 1.5260 2.5330 1.5760 ;
      RECT 2.4830 1.4280 2.5330 1.5260 ;
      RECT 2.4830 1.3780 3.2930 1.4280 ;
      RECT 3.2430 1.4280 3.2930 1.5440 ;
      RECT 4.5610 0.7360 4.9810 0.7860 ;
      RECT 4.5610 0.7860 4.6110 1.0990 ;
      RECT 4.0510 1.0990 4.6110 1.1490 ;
      RECT 4.0510 1.1490 4.1010 1.2720 ;
      RECT 3.8750 1.2720 4.1010 1.3220 ;
      RECT 3.8750 1.3220 3.9250 1.4280 ;
      RECT 3.6830 1.4280 3.9250 1.4780 ;
      RECT 4.5190 1.2080 4.9050 1.2580 ;
      RECT 3.3020 1.1660 3.6730 1.2160 ;
      RECT 3.6230 1.2160 3.6730 1.3080 ;
      RECT 3.6230 1.3080 3.8250 1.3580 ;
      RECT 3.7750 1.0510 3.8250 1.3080 ;
      RECT 3.7750 1.0060 3.8650 1.0510 ;
      RECT 2.7660 0.9560 3.8650 1.0060 ;
      RECT 3.8150 0.6560 3.8650 0.9560 ;
      RECT 3.7750 0.6060 3.8650 0.6560 ;
      RECT 3.7750 0.4960 3.8250 0.6060 ;
      RECT 3.6230 0.4460 3.8250 0.4960 ;
      RECT 3.6230 0.3710 3.6730 0.4460 ;
      RECT 3.7750 0.3710 3.8250 0.4460 ;
      RECT 2.6950 1.2780 3.0810 1.3280 ;
      RECT 4.4230 0.6340 5.5890 0.6840 ;
      RECT 4.4230 0.6840 4.4730 0.9780 ;
      RECT 4.0620 0.9780 4.4730 1.0280 ;
      RECT 4.0620 0.4960 4.1120 0.9780 ;
      RECT 4.0620 0.4460 4.1690 0.4960 ;
      RECT 4.4420 1.4080 4.9810 1.4580 ;
      RECT 2.6350 1.4780 3.1570 1.5280 ;
      RECT 2.6350 1.5280 2.6850 1.5650 ;
      RECT 0.8870 0.3120 1.5450 0.3620 ;
      RECT 0.8870 0.3620 0.9370 0.3940 ;
      RECT 1.4950 0.3620 1.5450 0.3940 ;
      RECT 1.7990 0.6180 2.2450 0.6680 ;
      RECT 1.7990 0.6680 1.8490 0.9140 ;
      RECT 1.7990 0.4220 1.8490 0.6180 ;
      RECT 2.2550 0.5180 2.3810 0.5680 ;
      RECT 2.2550 0.3940 2.3050 0.5180 ;
      RECT 2.3310 0.5680 2.3810 0.7180 ;
      RECT 2.2550 0.7180 2.3810 0.7680 ;
      RECT 2.2550 0.7680 2.3050 0.9140 ;
      RECT 0.7350 1.0420 0.9370 1.0920 ;
      RECT 0.8870 1.0920 0.9370 1.2160 ;
      RECT 0.7350 1.0920 0.7850 1.2160 ;
      RECT 0.7190 0.5120 1.2570 0.5620 ;
      RECT 2.0110 0.0960 2.7070 0.1460 ;
      RECT 1.1750 1.0880 1.5610 1.1380 ;
      RECT 1.4520 0.6040 1.6370 0.6540 ;
      RECT 0.2050 0.5280 0.2550 0.8880 ;
      RECT 0.2790 0.9380 0.3290 1.2160 ;
      RECT 0.2050 0.4780 0.3290 0.5280 ;
      RECT 0.2790 0.3180 0.3290 0.4780 ;
      RECT 0.2050 0.8880 1.5020 0.9380 ;
      RECT 1.4520 0.6540 1.5020 0.8880 ;
      RECT 4.4590 0.0880 4.5090 0.2300 ;
      RECT 3.5110 0.2300 4.5090 0.2800 ;
      RECT 3.8350 0.2800 3.9170 0.2900 ;
      RECT 3.5110 0.2800 3.5610 0.6040 ;
      RECT 3.0750 0.6040 3.5610 0.6540 ;
      RECT 3.8350 0.1880 3.9170 0.2300 ;
      RECT 2.5590 0.7560 3.4610 0.8060 ;
      RECT 2.5590 0.8060 2.6090 1.1580 ;
      RECT 2.5590 0.4840 2.6090 0.7560 ;
      RECT 2.5590 1.2080 2.6090 1.3140 ;
      RECT 2.5590 0.3550 2.6090 0.4340 ;
      RECT 2.5590 1.1580 2.9290 1.2080 ;
      RECT 2.5590 0.4340 2.7770 0.4840 ;
  END
END SDFFASRSX2_LVT

MACRO SDFFASRX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.08 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2950 0.8040 5.8410 0.8540 ;
        RECT 5.2950 0.8540 5.3450 1.5540 ;
        RECT 5.7910 0.5110 5.8410 0.8040 ;
        RECT 5.7210 0.4440 5.8410 0.5110 ;
        RECT 5.2950 0.3940 5.8410 0.4440 ;
        RECT 5.2950 0.1480 5.3450 0.3940 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 6.0800 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 1.6470 1.1340 1.6970 1.6420 ;
        RECT 5.1430 0.9120 5.1930 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 5.7510 1.0520 5.8010 1.6420 ;
        RECT 2.1030 1.3540 2.1530 1.6420 ;
        RECT 5.0310 1.3580 5.0810 1.6420 ;
        RECT 3.3430 1.3280 3.3930 1.6420 ;
        RECT 1.9510 1.3040 2.1530 1.3540 ;
        RECT 4.2020 1.3080 5.0810 1.3580 ;
        RECT 3.1500 1.2780 3.5520 1.3280 ;
        RECT 1.9510 1.0880 2.0010 1.3040 ;
        RECT 2.1030 1.1010 2.1530 1.3040 ;
    END
  END VDD

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8730 0.0970 5.9830 0.2070 ;
        RECT 5.9150 0.2070 5.9650 0.2700 ;
        RECT 5.5990 0.2700 5.9650 0.3200 ;
        RECT 5.5990 0.1480 5.6490 0.2700 ;
        RECT 5.9150 0.3200 5.9650 0.9180 ;
        RECT 5.5990 0.9180 5.9650 0.9680 ;
        RECT 5.5990 0.9680 5.6490 1.5460 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 0.6640 1.0110 0.8150 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END D

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9390 0.1060 4.2210 0.1560 ;
        RECT 4.1390 0.1560 4.2210 0.1920 ;
        RECT 2.9390 0.0970 3.0950 0.1060 ;
        RECT 2.9390 0.1560 3.0950 0.2350 ;
    END
    ANTENNAGATEAREA 0.0441 ;
  END RSTB

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6800 0.7250 0.7300 ;
        RECT 0.4010 0.5530 0.5110 0.6800 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2360 1.3150 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.7470 0.8570 4.9190 1.0340 ;
    END
    ANTENNAGATEAREA 0.0471 ;
  END SETB

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 6.0800 0.0300 ;
        RECT 1.6470 0.0300 1.6970 0.1960 ;
        RECT 5.1430 0.0300 5.1930 0.4080 ;
        RECT 0.5830 0.0300 0.6330 0.5150 ;
        RECT 5.7510 0.0300 5.8010 0.2200 ;
        RECT 0.4310 0.0300 0.4810 0.4370 ;
        RECT 2.7570 0.0300 2.8070 0.2870 ;
        RECT 4.9910 0.0300 5.0410 0.3580 ;
        RECT 1.6470 0.1960 2.1530 0.2460 ;
        RECT 2.7570 0.2870 3.3690 0.3370 ;
        RECT 4.3670 0.3580 5.0570 0.4080 ;
        RECT 2.1030 0.2460 2.1530 0.4500 ;
        RECT 1.9510 0.2460 2.0010 0.4500 ;
        RECT 1.6470 0.2460 1.6970 0.4080 ;
        RECT 3.3190 0.3370 3.3690 0.4610 ;
        RECT 3.1670 0.3370 3.2170 0.4610 ;
    END
  END VSS

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7690 1.4240 1.9410 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  OBS
    LAYER PO ;
      RECT 5.2290 0.0680 5.2590 1.6150 ;
      RECT 4.9250 0.9120 4.9550 1.6060 ;
      RECT 3.8610 0.0680 3.8910 0.6740 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 3.1010 0.7580 3.1310 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 5.0770 0.0680 5.1070 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 4.3170 0.0680 4.3470 1.6060 ;
      RECT 4.7730 0.0680 4.8030 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 3.7090 0.0680 3.7390 1.6060 ;
      RECT 4.4690 0.0680 4.4990 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 4.6210 0.0680 4.6510 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 2.4930 0.0680 2.5230 0.5920 ;
      RECT 2.4930 0.9900 2.5230 1.6060 ;
      RECT 4.9250 0.0680 4.9550 0.7870 ;
      RECT 3.1010 0.0680 3.1310 0.6290 ;
      RECT 3.8610 0.8820 3.8910 1.6060 ;
      RECT 5.8370 0.0680 5.8670 1.6060 ;
      RECT 5.6850 0.0680 5.7150 1.6060 ;
      RECT 5.9890 0.0680 6.0190 1.6060 ;
      RECT 5.5330 0.0680 5.5630 1.6060 ;
      RECT 5.3810 0.0680 5.4110 1.6060 ;
    LAYER NWELL ;
      RECT -0.1150 0.6790 6.1950 1.7730 ;
    LAYER M1 ;
      RECT 2.4070 1.0380 2.4570 1.3140 ;
      RECT 2.4310 0.3810 2.4810 0.9880 ;
      RECT 2.4070 0.2990 2.4970 0.3810 ;
      RECT 1.0230 0.9880 2.4810 1.0380 ;
      RECT 1.3430 0.4620 1.3930 0.5040 ;
      RECT 1.0230 0.4120 1.3930 0.4620 ;
      RECT 1.6870 0.5540 1.7370 0.7260 ;
      RECT 1.6500 0.7260 1.7370 0.7760 ;
      RECT 1.3430 0.5040 1.7370 0.5540 ;
      RECT 1.6500 0.7760 1.7000 0.9880 ;
      RECT 3.0750 0.7860 3.7650 0.8360 ;
      RECT 5.3800 0.6040 5.7410 0.6540 ;
      RECT 5.0310 0.7540 5.0810 1.1080 ;
      RECT 4.6710 1.1080 5.0810 1.1580 ;
      RECT 3.9270 0.4580 4.7540 0.5030 ;
      RECT 5.3800 0.6540 5.4300 0.7040 ;
      RECT 5.3800 0.5530 5.4300 0.6040 ;
      RECT 4.7040 0.5080 5.4300 0.5530 ;
      RECT 3.9270 0.5030 5.4300 0.5080 ;
      RECT 5.0310 0.7040 5.4300 0.7540 ;
      RECT 3.9270 0.5080 3.9770 1.1650 ;
      RECT 4.2300 0.5080 4.2800 0.7660 ;
      RECT 4.2300 0.7660 4.3730 0.8160 ;
      RECT 1.1750 1.0880 1.5610 1.1380 ;
      RECT 0.7350 1.0420 0.9370 1.0920 ;
      RECT 0.8870 1.0920 0.9370 1.2160 ;
      RECT 0.7350 1.0920 0.7850 1.2160 ;
      RECT 0.8870 0.3120 1.5450 0.3620 ;
      RECT 0.8870 0.3620 0.9370 0.3940 ;
      RECT 1.4950 0.3620 1.5450 0.3940 ;
      RECT 3.5020 1.5280 4.8420 1.5780 ;
      RECT 2.3150 1.5260 2.5330 1.5760 ;
      RECT 2.4830 1.4280 2.5330 1.5260 ;
      RECT 2.4830 1.3780 3.2930 1.4280 ;
      RECT 3.2430 1.4280 3.2930 1.5440 ;
      RECT 4.5610 0.7090 4.9810 0.7590 ;
      RECT 4.5610 0.7590 4.6110 1.0990 ;
      RECT 4.0510 1.0990 4.6110 1.1490 ;
      RECT 4.0510 1.1490 4.1010 1.2720 ;
      RECT 3.8750 1.2720 4.1010 1.3220 ;
      RECT 3.8750 1.3220 3.9250 1.4280 ;
      RECT 3.6830 1.4280 3.9250 1.4780 ;
      RECT 4.5190 1.2080 4.9050 1.2580 ;
      RECT 3.3020 1.1660 3.6730 1.2160 ;
      RECT 3.6230 1.2160 3.6730 1.3080 ;
      RECT 3.6230 1.3080 3.8250 1.3580 ;
      RECT 3.7750 1.0510 3.8250 1.3080 ;
      RECT 2.7660 1.0010 3.8650 1.0510 ;
      RECT 3.8150 0.6560 3.8650 1.0010 ;
      RECT 3.7750 0.6060 3.8650 0.6560 ;
      RECT 3.7750 0.4960 3.8250 0.6060 ;
      RECT 3.6230 0.4460 3.8250 0.4960 ;
      RECT 3.6230 0.3710 3.6730 0.4460 ;
      RECT 3.7750 0.3710 3.8250 0.4460 ;
      RECT 2.6950 1.2780 3.0810 1.3280 ;
      RECT 4.4230 0.6040 5.3140 0.6540 ;
      RECT 4.4230 0.6540 4.4730 0.9780 ;
      RECT 4.0620 0.9780 4.4730 1.0280 ;
      RECT 4.0620 0.6080 4.1120 0.9780 ;
      RECT 4.0620 0.5580 4.1690 0.6080 ;
      RECT 4.4420 1.4080 4.9810 1.4580 ;
      RECT 2.6350 1.4780 3.1570 1.5280 ;
      RECT 2.6350 1.5280 2.6850 1.5650 ;
      RECT 1.7990 0.6180 2.2450 0.6680 ;
      RECT 1.7990 0.6680 1.8490 0.9140 ;
      RECT 1.7990 0.4220 1.8490 0.6180 ;
      RECT 2.2550 0.5180 2.3810 0.5680 ;
      RECT 2.2550 0.3940 2.3050 0.5180 ;
      RECT 2.3310 0.5680 2.3810 0.7180 ;
      RECT 2.2550 0.7180 2.3810 0.7680 ;
      RECT 2.2550 0.7680 2.3050 0.9140 ;
      RECT 0.7190 0.5120 1.2570 0.5620 ;
      RECT 2.0110 0.0960 2.7070 0.1460 ;
      RECT 1.4520 0.6040 1.6370 0.6540 ;
      RECT 0.2050 0.5280 0.2550 0.8880 ;
      RECT 0.2790 0.9380 0.3290 1.2160 ;
      RECT 0.2050 0.4780 0.3290 0.5280 ;
      RECT 0.2790 0.3180 0.3290 0.4780 ;
      RECT 0.2050 0.8880 1.5020 0.9380 ;
      RECT 1.4520 0.6540 1.5020 0.8880 ;
      RECT 4.4590 0.1520 4.5090 0.2580 ;
      RECT 3.5110 0.2580 4.5090 0.3080 ;
      RECT 3.5110 0.2300 3.5610 0.2580 ;
      RECT 3.5110 0.3080 3.5610 0.5720 ;
      RECT 3.0750 0.5720 3.5610 0.6220 ;
      RECT 3.8350 0.2060 3.9170 0.2580 ;
      RECT 2.5590 0.6720 3.4610 0.7220 ;
      RECT 2.5590 0.7220 2.6090 1.1580 ;
      RECT 2.5590 0.4840 2.6090 0.6720 ;
      RECT 2.5590 1.2080 2.6090 1.3140 ;
      RECT 2.5590 0.3550 2.6090 0.4340 ;
      RECT 2.5590 1.1580 2.9290 1.2080 ;
      RECT 2.5590 0.4340 2.7770 0.4840 ;
  END
END SDFFASRX1_LVT

MACRO SDFFASRX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.08 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2950 0.8040 5.8410 0.8540 ;
        RECT 5.2950 0.8540 5.3450 1.5460 ;
        RECT 5.7910 0.5110 5.8410 0.8040 ;
        RECT 5.7210 0.4440 5.8410 0.5110 ;
        RECT 5.2950 0.3940 5.8410 0.4440 ;
        RECT 5.2950 0.1480 5.3450 0.3940 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 6.0800 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 5.4470 0.9600 5.4970 1.6420 ;
        RECT 1.6470 1.1340 1.6970 1.6420 ;
        RECT 5.1430 0.9120 5.1930 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 5.7510 1.0520 5.8010 1.6420 ;
        RECT 3.3430 1.3280 3.3930 1.6420 ;
        RECT 2.1030 1.3540 2.1530 1.6420 ;
        RECT 5.0310 1.3580 5.0810 1.6420 ;
        RECT 3.1500 1.2780 3.5520 1.3280 ;
        RECT 1.9510 1.3040 2.1530 1.3540 ;
        RECT 4.2020 1.3080 5.0810 1.3580 ;
        RECT 1.9510 1.0880 2.0010 1.3040 ;
        RECT 2.1030 1.1010 2.1530 1.3040 ;
    END
  END VDD

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8730 0.0970 5.9830 0.2070 ;
        RECT 5.9150 0.2070 5.9650 0.2700 ;
        RECT 5.5990 0.2700 5.9650 0.3200 ;
        RECT 5.5990 0.1480 5.6490 0.2700 ;
        RECT 5.9150 0.3200 5.9650 0.9180 ;
        RECT 5.5990 0.9180 5.9650 0.9680 ;
        RECT 5.5990 0.9680 5.6490 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 0.6640 1.0110 0.8150 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END D

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9390 0.0880 4.2210 0.1380 ;
        RECT 4.1390 0.1380 4.2210 0.1740 ;
        RECT 2.9390 0.1380 3.0950 0.2070 ;
    END
    ANTENNAGATEAREA 0.0441 ;
  END RSTB

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6800 0.7250 0.7300 ;
        RECT 0.4010 0.5530 0.5110 0.6800 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2360 1.3150 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.7470 0.8570 4.9190 1.0340 ;
    END
    ANTENNAGATEAREA 0.0471 ;
  END SETB

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 6.0800 0.0300 ;
        RECT 1.6470 0.0300 1.6970 0.1960 ;
        RECT 5.1430 0.0300 5.1930 0.4080 ;
        RECT 5.4470 0.0300 5.4970 0.3190 ;
        RECT 0.5830 0.0300 0.6330 0.5150 ;
        RECT 5.7510 0.0300 5.8010 0.2200 ;
        RECT 0.4310 0.0300 0.4810 0.4370 ;
        RECT 2.7570 0.0300 2.8070 0.2870 ;
        RECT 4.9910 0.0300 5.0410 0.3300 ;
        RECT 1.6470 0.1960 2.1530 0.2460 ;
        RECT 2.7570 0.2870 3.3690 0.3370 ;
        RECT 4.3670 0.3300 5.0570 0.3800 ;
        RECT 2.1030 0.2460 2.1530 0.4500 ;
        RECT 1.9510 0.2460 2.0010 0.4500 ;
        RECT 1.6470 0.2460 1.6970 0.4080 ;
        RECT 3.3190 0.3370 3.3690 0.4610 ;
        RECT 3.1670 0.3370 3.2170 0.4610 ;
    END
  END VSS

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7690 1.4240 1.9410 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  OBS
    LAYER PO ;
      RECT 5.5330 0.0680 5.5630 1.6060 ;
      RECT 5.3810 0.0680 5.4110 1.6060 ;
      RECT 5.2290 0.0680 5.2590 1.6060 ;
      RECT 4.9250 0.9120 4.9550 1.6060 ;
      RECT 3.8610 0.0680 3.8910 0.6320 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 3.1010 0.7580 3.1310 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 5.0770 0.0680 5.1070 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 4.3170 0.0680 4.3470 1.6060 ;
      RECT 4.7730 0.0680 4.8030 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 3.7090 0.0680 3.7390 1.6060 ;
      RECT 4.4690 0.0680 4.4990 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 4.6210 0.0680 4.6510 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 2.4930 0.0680 2.5230 0.5920 ;
      RECT 2.4930 0.9900 2.5230 1.6060 ;
      RECT 4.9250 0.0680 4.9550 0.7870 ;
      RECT 3.1010 0.0680 3.1310 0.6180 ;
      RECT 3.8610 0.8820 3.8910 1.6060 ;
      RECT 5.8370 0.0680 5.8670 1.6060 ;
      RECT 5.6850 0.0680 5.7150 1.6060 ;
      RECT 5.9890 0.0680 6.0190 1.6060 ;
    LAYER NWELL ;
      RECT -0.1150 0.6790 6.1950 1.7730 ;
    LAYER M1 ;
      RECT 2.4070 1.0380 2.4570 1.3140 ;
      RECT 2.4310 0.3810 2.4810 0.9880 ;
      RECT 2.4070 0.2990 2.4970 0.3810 ;
      RECT 1.0230 0.9880 2.4810 1.0380 ;
      RECT 1.3430 0.4620 1.3930 0.5040 ;
      RECT 1.0230 0.4120 1.3930 0.4620 ;
      RECT 1.6500 0.7760 1.7000 0.9880 ;
      RECT 1.6500 0.7260 1.7370 0.7760 ;
      RECT 1.6870 0.5540 1.7370 0.7260 ;
      RECT 1.3430 0.5040 1.7370 0.5540 ;
      RECT 3.0750 0.7860 3.7650 0.8360 ;
      RECT 5.5040 0.6040 5.7410 0.6540 ;
      RECT 5.5040 0.6540 5.5540 0.7040 ;
      RECT 5.5040 0.5530 5.5540 0.6040 ;
      RECT 4.7040 0.5030 5.5540 0.5530 ;
      RECT 5.0310 0.7040 5.5540 0.7540 ;
      RECT 5.0310 0.7540 5.0810 1.1080 ;
      RECT 4.7040 0.4880 4.7540 0.5030 ;
      RECT 4.6710 1.1080 5.0810 1.1580 ;
      RECT 3.9270 0.4380 4.7540 0.4880 ;
      RECT 3.9270 0.4880 3.9770 1.1650 ;
      RECT 4.2300 0.4880 4.2800 0.7660 ;
      RECT 4.2300 0.7660 4.3730 0.8160 ;
      RECT 1.1750 1.0880 1.5610 1.1380 ;
      RECT 0.7350 1.0420 0.9370 1.0920 ;
      RECT 0.8870 1.0920 0.9370 1.2160 ;
      RECT 0.7350 1.0920 0.7850 1.2160 ;
      RECT 0.8870 0.3120 1.5450 0.3620 ;
      RECT 0.8870 0.3620 0.9370 0.3940 ;
      RECT 1.4950 0.3620 1.5450 0.3940 ;
      RECT 3.5020 1.5280 4.8420 1.5780 ;
      RECT 2.3150 1.5260 2.5330 1.5760 ;
      RECT 2.4830 1.4280 2.5330 1.5260 ;
      RECT 2.4830 1.3780 3.2930 1.4280 ;
      RECT 3.2430 1.4280 3.2930 1.5440 ;
      RECT 4.5610 0.7090 4.9810 0.7590 ;
      RECT 4.5610 0.7590 4.6110 1.0990 ;
      RECT 4.0510 1.0990 4.6110 1.1490 ;
      RECT 4.0510 1.1490 4.1010 1.2720 ;
      RECT 3.8750 1.2720 4.1010 1.3220 ;
      RECT 3.8750 1.3220 3.9250 1.4280 ;
      RECT 3.6830 1.4280 3.9250 1.4780 ;
      RECT 4.5190 1.2080 4.9050 1.2580 ;
      RECT 3.3020 1.1660 3.6730 1.2160 ;
      RECT 3.6230 1.2160 3.6730 1.3080 ;
      RECT 3.6230 1.3080 3.8250 1.3580 ;
      RECT 3.7750 1.0510 3.8250 1.3080 ;
      RECT 2.7660 1.0010 3.8650 1.0510 ;
      RECT 3.8150 0.6560 3.8650 1.0010 ;
      RECT 3.7750 0.6060 3.8650 0.6560 ;
      RECT 3.7750 0.4960 3.8250 0.6060 ;
      RECT 3.6230 0.4460 3.8250 0.4960 ;
      RECT 3.6230 0.3710 3.6730 0.4460 ;
      RECT 3.7750 0.3710 3.8250 0.4460 ;
      RECT 2.6950 1.2780 3.0810 1.3280 ;
      RECT 4.4230 0.6040 5.4370 0.6540 ;
      RECT 4.4230 0.6540 4.4730 0.9780 ;
      RECT 4.0620 0.9780 4.4730 1.0280 ;
      RECT 4.0620 0.5880 4.1120 0.9780 ;
      RECT 4.0620 0.5380 4.1690 0.5880 ;
      RECT 4.4420 1.4080 4.9810 1.4580 ;
      RECT 2.6350 1.4780 3.1570 1.5280 ;
      RECT 2.6350 1.5280 2.6850 1.5650 ;
      RECT 1.7990 0.6180 2.2450 0.6680 ;
      RECT 1.7990 0.6680 1.8490 0.9140 ;
      RECT 1.7990 0.4220 1.8490 0.6180 ;
      RECT 2.2550 0.5180 2.3810 0.5680 ;
      RECT 2.2550 0.3940 2.3050 0.5180 ;
      RECT 2.3310 0.5680 2.3810 0.7180 ;
      RECT 2.2550 0.7180 2.3810 0.7680 ;
      RECT 2.2550 0.7680 2.3050 0.9140 ;
      RECT 0.7190 0.5120 1.2570 0.5620 ;
      RECT 2.0110 0.0960 2.7070 0.1460 ;
      RECT 1.4520 0.6040 1.6370 0.6540 ;
      RECT 0.2050 0.5280 0.2550 0.8880 ;
      RECT 0.2790 0.9380 0.3290 1.2160 ;
      RECT 0.2050 0.4780 0.3290 0.5280 ;
      RECT 0.2790 0.3180 0.3290 0.4780 ;
      RECT 0.2050 0.8880 1.5020 0.9380 ;
      RECT 1.4520 0.6540 1.5020 0.8880 ;
      RECT 4.4590 0.0880 4.5090 0.2300 ;
      RECT 3.5110 0.2300 4.5090 0.2800 ;
      RECT 3.8350 0.2800 3.9170 0.2900 ;
      RECT 3.5110 0.2800 3.5610 0.5400 ;
      RECT 3.0750 0.5400 3.5610 0.5900 ;
      RECT 3.8350 0.1880 3.9170 0.2300 ;
      RECT 2.5590 0.6400 3.4610 0.6900 ;
      RECT 2.5590 0.6900 2.6090 1.1580 ;
      RECT 2.5590 0.4840 2.6090 0.6400 ;
      RECT 2.5590 1.2080 2.6090 1.3140 ;
      RECT 2.5590 0.3550 2.6090 0.4340 ;
      RECT 2.5590 1.1580 2.9290 1.2080 ;
      RECT 2.5590 0.4340 2.7770 0.4840 ;
  END
END SDFFASRX2_LVT

MACRO SDFFASX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.472 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2360 1.3150 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4430 0.8570 4.6150 1.0340 ;
    END
    ANTENNAGATEAREA 0.0441 ;
  END SETB

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2650 1.1610 5.3760 1.2210 ;
        RECT 5.1430 1.2210 5.3760 1.2710 ;
        RECT 5.3250 0.2040 5.3750 1.1610 ;
        RECT 5.1430 1.2710 5.1930 1.5460 ;
        RECT 5.1270 0.1540 5.3750 0.2040 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6800 0.7250 0.7300 ;
        RECT 0.4010 0.5530 0.5110 0.6800 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 0.6640 1.0110 0.8150 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 5.4720 0.0300 ;
        RECT 1.8020 0.0300 1.8520 0.1960 ;
        RECT 0.4310 0.0300 0.4810 0.4370 ;
        RECT 0.5830 0.0300 0.6330 0.5150 ;
        RECT 1.6470 0.0300 1.6970 0.4080 ;
        RECT 3.1670 0.0300 3.2170 0.4610 ;
        RECT 4.9910 0.0300 5.0410 0.2200 ;
        RECT 3.0150 0.0300 3.0650 0.3710 ;
        RECT 4.6870 0.0300 4.7370 0.3350 ;
        RECT 1.8020 0.1960 2.1530 0.2460 ;
        RECT 4.0610 0.3350 4.7530 0.3850 ;
        RECT 1.9510 0.2460 2.0010 0.4500 ;
        RECT 2.1030 0.2460 2.1530 0.4500 ;
    END
  END VSS

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.1130 1.0090 5.2230 1.1190 ;
        RECT 5.1730 0.8540 5.2230 1.0090 ;
        RECT 4.8390 0.8040 5.2230 0.8540 ;
        RECT 4.8390 0.8540 4.8890 1.5460 ;
        RECT 5.1730 0.3590 5.2230 0.8040 ;
        RECT 4.8390 0.3090 5.2230 0.3590 ;
        RECT 4.8390 0.1480 4.8890 0.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7690 1.4240 1.9410 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 5.4720 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 4.9910 0.9470 5.0410 1.6420 ;
        RECT 2.1030 1.3540 2.1530 1.6420 ;
        RECT 3.1910 1.3210 3.2410 1.6420 ;
        RECT 4.7270 1.3580 4.7770 1.6420 ;
        RECT 1.6470 1.3400 1.6990 1.6420 ;
        RECT 1.9510 1.3040 2.1530 1.3540 ;
        RECT 2.9900 1.2710 3.4000 1.3210 ;
        RECT 4.0500 1.3080 4.7770 1.3580 ;
        RECT 1.6470 1.1340 1.6970 1.3400 ;
        RECT 1.9510 1.0880 2.0010 1.3040 ;
        RECT 2.1030 1.1010 2.1530 1.3040 ;
    END
  END VDD
  OBS
    LAYER PO ;
      RECT 2.9490 0.7280 2.9790 1.6040 ;
      RECT 2.6450 0.0660 2.6750 1.6040 ;
      RECT 4.6210 1.0120 4.6510 1.6060 ;
      RECT 4.6210 0.0680 4.6510 0.7870 ;
      RECT 3.7090 0.8820 3.7390 1.6060 ;
      RECT 4.0130 0.0650 4.0430 1.6030 ;
      RECT 5.3810 0.0680 5.4110 1.6060 ;
      RECT 4.9250 0.0680 4.9550 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6040 ;
      RECT 3.1010 0.0660 3.1310 1.6040 ;
      RECT 4.3170 0.0680 4.3470 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 5.0770 0.0680 5.1070 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 4.4690 0.0680 4.4990 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 5.2290 0.0680 5.2590 1.6060 ;
      RECT 4.7730 0.0680 4.8030 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 2.4930 0.0680 2.5230 0.5420 ;
      RECT 2.9490 0.0660 2.9790 0.6160 ;
      RECT 2.4930 0.9900 2.5230 1.6060 ;
      RECT 3.7090 0.0680 3.7390 0.6220 ;
    LAYER NWELL ;
      RECT 3.8760 0.6690 4.1800 0.6790 ;
      RECT -0.1150 0.6790 5.5870 1.7730 ;
    LAYER M1 ;
      RECT 3.0910 1.4260 3.1410 1.5600 ;
      RECT 2.4830 1.3760 3.1410 1.4260 ;
      RECT 2.4830 1.4260 2.5330 1.5260 ;
      RECT 2.3150 1.5260 2.5330 1.5760 ;
      RECT 3.6230 0.6060 3.7130 0.6560 ;
      RECT 3.6630 0.6560 3.7130 1.0010 ;
      RECT 3.6230 0.4960 3.6730 0.6060 ;
      RECT 2.7660 1.0010 3.7130 1.0510 ;
      RECT 3.4710 0.4460 3.6730 0.4960 ;
      RECT 3.6230 1.0510 3.6730 1.3080 ;
      RECT 3.4710 0.3710 3.5210 0.4460 ;
      RECT 3.6230 0.3710 3.6730 0.4460 ;
      RECT 3.4710 1.3080 3.6730 1.3580 ;
      RECT 3.4710 1.2160 3.5210 1.3080 ;
      RECT 3.1500 1.1660 3.5210 1.2160 ;
      RECT 2.6350 1.4760 3.0050 1.5260 ;
      RECT 2.6350 1.5260 2.6850 1.5630 ;
      RECT 4.1480 0.6040 4.9810 0.6540 ;
      RECT 4.1480 0.6540 4.1980 0.9750 ;
      RECT 4.1480 0.5850 4.1980 0.6040 ;
      RECT 3.9040 0.9750 4.1980 1.0250 ;
      RECT 3.9110 0.5350 4.1980 0.5850 ;
      RECT 3.3500 1.5170 3.8980 1.5670 ;
      RECT 3.8480 1.4610 3.8980 1.5170 ;
      RECT 3.8480 1.4110 4.5250 1.4610 ;
      RECT 0.7350 1.0420 0.9370 1.0920 ;
      RECT 0.7350 1.0920 0.7850 1.2160 ;
      RECT 0.8870 1.0920 0.9370 1.2160 ;
      RECT 0.8870 0.3120 1.5450 0.3620 ;
      RECT 1.4950 0.3620 1.5450 0.3940 ;
      RECT 0.8870 0.3620 0.9370 0.3940 ;
      RECT 0.7190 0.5120 1.2570 0.5620 ;
      RECT 4.2670 0.7090 4.6770 0.7590 ;
      RECT 4.2670 0.7590 4.3170 1.0990 ;
      RECT 3.8990 1.0990 4.3170 1.1490 ;
      RECT 3.8990 1.1490 3.9490 1.2720 ;
      RECT 3.8990 1.0960 3.9490 1.0990 ;
      RECT 3.7230 1.2720 3.9490 1.3220 ;
      RECT 3.7230 1.3220 3.7730 1.4170 ;
      RECT 3.5310 1.4170 3.7730 1.4670 ;
      RECT 2.2550 0.5180 2.3810 0.5680 ;
      RECT 2.2550 0.3940 2.3050 0.5180 ;
      RECT 2.3310 0.5680 2.3810 0.7180 ;
      RECT 2.2550 0.7180 2.3810 0.7680 ;
      RECT 2.2550 0.7680 2.3050 0.9140 ;
      RECT 1.1750 1.0880 1.5610 1.1380 ;
      RECT 4.2150 1.2080 4.6010 1.2580 ;
      RECT 4.1380 1.5280 4.6770 1.5780 ;
      RECT 1.7990 0.6180 2.2450 0.6680 ;
      RECT 1.7990 0.6680 1.8490 0.9140 ;
      RECT 1.7990 0.4220 1.8490 0.6180 ;
      RECT 2.0110 0.0960 2.7070 0.1460 ;
      RECT 3.3590 0.2300 4.2050 0.2800 ;
      RECT 4.1550 0.1330 4.2050 0.2300 ;
      RECT 3.6830 0.1780 3.7650 0.2300 ;
      RECT 3.3590 0.2800 3.4090 0.5380 ;
      RECT 2.9220 0.5380 3.4090 0.5880 ;
      RECT 3.3590 0.5880 3.4090 0.5900 ;
      RECT 2.9140 0.7560 3.6130 0.8060 ;
      RECT 2.4070 0.2990 2.4970 0.3810 ;
      RECT 2.4310 0.3810 2.4810 0.9880 ;
      RECT 2.4070 1.0380 2.4570 1.3140 ;
      RECT 1.0230 0.9880 2.4810 1.0380 ;
      RECT 1.3430 0.4620 1.3930 0.5040 ;
      RECT 1.0230 0.4120 1.3930 0.4620 ;
      RECT 1.6500 0.7760 1.7000 0.9880 ;
      RECT 1.6500 0.7260 1.7370 0.7760 ;
      RECT 1.6870 0.5540 1.7370 0.7260 ;
      RECT 1.3430 0.5040 1.7370 0.5540 ;
      RECT 5.0670 0.4850 5.1170 0.7040 ;
      RECT 3.7750 0.4350 5.1170 0.4850 ;
      RECT 4.7270 0.7040 5.1170 0.7540 ;
      RECT 4.7270 0.7540 4.7770 1.1080 ;
      RECT 4.3670 1.1080 4.7770 1.1580 ;
      RECT 3.7750 0.4850 3.8250 0.6350 ;
      RECT 3.7750 0.6350 4.0690 0.6850 ;
      RECT 3.7750 0.6850 3.8250 1.1650 ;
      RECT 2.5590 0.6400 3.3090 0.6900 ;
      RECT 2.5590 0.6900 2.6090 1.1560 ;
      RECT 2.5590 0.4820 2.6090 0.6400 ;
      RECT 2.5590 1.1560 2.7770 1.2060 ;
      RECT 2.5590 0.4320 2.7770 0.4820 ;
      RECT 2.5590 1.2060 2.6090 1.3140 ;
      RECT 2.5590 0.3550 2.6090 0.4320 ;
      RECT 1.4520 0.6040 1.6370 0.6540 ;
      RECT 0.2050 0.5280 0.2550 0.8880 ;
      RECT 0.2790 0.9380 0.3290 1.2160 ;
      RECT 0.2050 0.4780 0.3290 0.5280 ;
      RECT 0.2790 0.3180 0.3290 0.4780 ;
      RECT 0.2050 0.8880 1.5020 0.9380 ;
      RECT 1.4520 0.6540 1.5020 0.8880 ;
  END
END SDFFASX1_LVT

MACRO SDFFASX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.776 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.9910 0.1480 5.0410 0.3940 ;
        RECT 4.9910 0.3940 5.5370 0.4440 ;
        RECT 5.4170 0.4440 5.5370 0.5110 ;
        RECT 5.4870 0.5110 5.5370 0.8040 ;
        RECT 4.9910 0.8040 5.5370 0.8540 ;
        RECT 4.9910 0.8540 5.0410 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.5690 0.0970 5.6790 0.2070 ;
        RECT 5.6110 0.2070 5.6610 0.2700 ;
        RECT 5.2950 0.2700 5.6610 0.3200 ;
        RECT 5.2950 0.1480 5.3450 0.2700 ;
        RECT 5.6110 0.3200 5.6610 0.9180 ;
        RECT 5.2950 0.9180 5.6610 0.9680 ;
        RECT 5.2950 0.9680 5.3450 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2360 1.3150 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4430 0.8570 4.6150 1.0340 ;
    END
    ANTENNAGATEAREA 0.0441 ;
  END SETB

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6800 0.7250 0.7300 ;
        RECT 0.4010 0.5530 0.5110 0.6800 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 0.6640 1.0110 0.8150 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 5.7760 0.0300 ;
        RECT 1.8020 0.0300 1.8520 0.1960 ;
        RECT 0.4310 0.0300 0.4810 0.4370 ;
        RECT 0.5830 0.0300 0.6330 0.5150 ;
        RECT 5.4470 0.0300 5.4970 0.2200 ;
        RECT 4.8390 0.0300 4.8890 0.4080 ;
        RECT 5.1430 0.0300 5.1930 0.3190 ;
        RECT 1.6470 0.0300 1.6970 0.4080 ;
        RECT 3.1670 0.0300 3.2170 0.4610 ;
        RECT 4.6870 0.0300 4.7370 0.3430 ;
        RECT 3.0150 0.0300 3.0650 0.3710 ;
        RECT 1.8020 0.1960 2.1530 0.2460 ;
        RECT 4.0610 0.3430 4.7530 0.3930 ;
        RECT 1.9510 0.2460 2.0010 0.4500 ;
        RECT 2.1030 0.2460 2.1530 0.4500 ;
    END
  END VSS

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7690 1.4240 1.9410 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 5.7760 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 5.4470 1.0520 5.4970 1.6420 ;
        RECT 5.1430 0.9600 5.1930 1.6420 ;
        RECT 4.8390 0.9120 4.8890 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 2.1030 1.3540 2.1530 1.6420 ;
        RECT 3.1910 1.3210 3.2410 1.6420 ;
        RECT 4.7270 1.3580 4.7770 1.6420 ;
        RECT 1.6470 1.3400 1.6990 1.6420 ;
        RECT 1.9510 1.3040 2.1530 1.3540 ;
        RECT 2.9900 1.2710 3.4000 1.3210 ;
        RECT 4.0500 1.3080 4.7770 1.3580 ;
        RECT 1.6470 1.1340 1.6970 1.3400 ;
        RECT 1.9510 1.0880 2.0010 1.3040 ;
        RECT 2.1030 1.1010 2.1530 1.3040 ;
    END
  END VDD
  OBS
    LAYER PO ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 5.5330 0.0680 5.5630 1.6060 ;
      RECT 5.3810 0.0680 5.4110 1.6060 ;
      RECT 5.6850 0.0680 5.7150 1.6060 ;
      RECT 5.2290 0.0680 5.2590 1.6060 ;
      RECT 5.0770 0.0680 5.1070 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 4.4690 0.0680 4.4990 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 4.7730 0.0680 4.8030 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 2.4930 0.0680 2.5230 0.5420 ;
      RECT 2.9490 0.0660 2.9790 0.6160 ;
      RECT 2.4930 0.9900 2.5230 1.6060 ;
      RECT 3.7090 0.0680 3.7390 0.6220 ;
      RECT 2.9490 0.7280 2.9790 1.6040 ;
      RECT 2.6450 0.0660 2.6750 1.6040 ;
      RECT 4.6210 1.0120 4.6510 1.6060 ;
      RECT 4.6210 0.0680 4.6510 0.7870 ;
      RECT 3.7090 0.8820 3.7390 1.6060 ;
      RECT 4.0130 0.0650 4.0430 1.6030 ;
      RECT 4.9250 0.0680 4.9550 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6040 ;
      RECT 3.1010 0.0660 3.1310 1.6040 ;
      RECT 4.3170 0.0680 4.3470 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
    LAYER NWELL ;
      RECT -0.1150 0.6790 5.8910 1.7730 ;
      RECT 3.8760 0.6750 4.1800 0.6790 ;
    LAYER M1 ;
      RECT 2.5590 0.6400 3.3090 0.6900 ;
      RECT 2.5590 1.2060 2.6090 1.3140 ;
      RECT 2.5590 1.1560 2.7770 1.2060 ;
      RECT 2.5590 0.6900 2.6090 1.1560 ;
      RECT 2.5590 0.4820 2.6090 0.6400 ;
      RECT 2.5590 0.4320 2.7770 0.4820 ;
      RECT 2.5590 0.3550 2.6090 0.4320 ;
      RECT 1.4520 0.6040 1.6370 0.6540 ;
      RECT 0.2050 0.5280 0.2550 0.8880 ;
      RECT 0.2790 0.9380 0.3290 1.2160 ;
      RECT 0.2050 0.4780 0.3290 0.5280 ;
      RECT 0.2790 0.3180 0.3290 0.4780 ;
      RECT 0.2050 0.8880 1.5020 0.9380 ;
      RECT 1.4520 0.6540 1.5020 0.8880 ;
      RECT 3.6230 0.6060 3.7130 0.6560 ;
      RECT 3.6230 0.4960 3.6730 0.6060 ;
      RECT 3.6630 0.6560 3.7130 1.0010 ;
      RECT 3.4710 0.4460 3.6730 0.4960 ;
      RECT 2.7660 1.0010 3.7130 1.0510 ;
      RECT 3.6230 0.3710 3.6730 0.4460 ;
      RECT 3.4710 0.3710 3.5210 0.4460 ;
      RECT 3.6230 1.0510 3.6730 1.3080 ;
      RECT 3.4710 1.3080 3.6730 1.3580 ;
      RECT 3.4710 1.2160 3.5210 1.3080 ;
      RECT 3.1500 1.1660 3.5210 1.2160 ;
      RECT 4.1480 0.6040 5.1330 0.6540 ;
      RECT 4.1480 0.6540 4.1980 0.9750 ;
      RECT 4.1480 0.5930 4.1980 0.6040 ;
      RECT 3.9110 0.9750 4.1980 1.0250 ;
      RECT 3.9110 0.5430 4.1980 0.5930 ;
      RECT 2.0110 0.0960 2.7070 0.1460 ;
      RECT 2.6350 1.4760 3.0050 1.5260 ;
      RECT 2.6350 1.5260 2.6850 1.5630 ;
      RECT 2.3150 1.5260 2.5330 1.5760 ;
      RECT 2.4830 1.4260 2.5330 1.5260 ;
      RECT 2.4830 1.3760 3.1410 1.4260 ;
      RECT 3.0910 1.4260 3.1410 1.5840 ;
      RECT 3.3500 1.5280 3.8980 1.5780 ;
      RECT 3.8480 1.4610 3.8980 1.5280 ;
      RECT 3.8480 1.4110 4.5250 1.4610 ;
      RECT 0.7350 1.0420 0.9370 1.0920 ;
      RECT 0.7350 1.0920 0.7850 1.2160 ;
      RECT 0.8870 1.0920 0.9370 1.2160 ;
      RECT 0.8870 0.3120 1.5450 0.3620 ;
      RECT 1.4950 0.3620 1.5450 0.3940 ;
      RECT 0.8870 0.3620 0.9370 0.3940 ;
      RECT 0.7190 0.5120 1.2570 0.5620 ;
      RECT 4.2670 0.7090 4.6770 0.7590 ;
      RECT 4.2670 0.7590 4.3170 1.0990 ;
      RECT 3.8990 1.0990 4.3170 1.1490 ;
      RECT 3.8990 1.1490 3.9490 1.2720 ;
      RECT 3.8990 1.0960 3.9490 1.0990 ;
      RECT 3.7230 1.2720 3.9490 1.3220 ;
      RECT 3.7230 1.3220 3.7730 1.4280 ;
      RECT 3.5310 1.4280 3.7730 1.4780 ;
      RECT 2.2550 0.5180 2.3810 0.5680 ;
      RECT 2.2550 0.3940 2.3050 0.5180 ;
      RECT 2.3310 0.5680 2.3810 0.7180 ;
      RECT 2.2550 0.7180 2.3810 0.7680 ;
      RECT 2.2550 0.7680 2.3050 0.9140 ;
      RECT 1.1750 1.0880 1.5610 1.1380 ;
      RECT 4.2150 1.2080 4.6010 1.2580 ;
      RECT 4.1380 1.5340 4.6770 1.5840 ;
      RECT 1.7990 0.6180 2.2450 0.6680 ;
      RECT 1.7990 0.6680 1.8490 0.9140 ;
      RECT 1.7990 0.4220 1.8490 0.6180 ;
      RECT 3.3590 0.1940 4.2050 0.2440 ;
      RECT 4.1550 0.0880 4.2050 0.1940 ;
      RECT 3.6830 0.1420 3.7650 0.1940 ;
      RECT 3.3590 0.2440 3.4090 0.5380 ;
      RECT 2.9220 0.5380 3.4090 0.5880 ;
      RECT 3.3590 0.5880 3.4090 0.5900 ;
      RECT 2.9140 0.7560 3.6130 0.8060 ;
      RECT 2.4070 0.2990 2.4970 0.3810 ;
      RECT 2.4310 0.3810 2.4810 0.9880 ;
      RECT 2.4070 1.0380 2.4570 1.3140 ;
      RECT 1.0230 0.9880 2.4810 1.0380 ;
      RECT 1.3430 0.4620 1.3930 0.5040 ;
      RECT 1.0230 0.4120 1.3930 0.4620 ;
      RECT 1.6500 0.7760 1.7000 0.9880 ;
      RECT 1.6500 0.7260 1.7370 0.7760 ;
      RECT 1.6870 0.5540 1.7370 0.7260 ;
      RECT 1.3430 0.5040 1.7370 0.5540 ;
      RECT 5.2000 0.6040 5.4370 0.6540 ;
      RECT 4.7270 0.7540 4.7770 1.1080 ;
      RECT 4.4240 0.4930 4.4740 0.5030 ;
      RECT 4.3670 1.1080 4.7770 1.1580 ;
      RECT 3.7750 0.4430 4.4740 0.4930 ;
      RECT 3.7750 0.4930 3.8250 0.6460 ;
      RECT 3.7750 0.6460 4.0690 0.6960 ;
      RECT 3.7750 0.6960 3.8250 1.1650 ;
      RECT 5.2000 0.6540 5.2500 0.7040 ;
      RECT 5.2000 0.5530 5.2500 0.6040 ;
      RECT 4.4240 0.5030 5.2500 0.5530 ;
      RECT 4.7270 0.7040 5.2500 0.7540 ;
  END
END SDFFASX2_LVT

MACRO SDFFNARX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.472 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 5.4720 0.0300 ;
        RECT 1.8020 0.0300 1.8520 0.1960 ;
        RECT 0.4310 0.0300 0.4810 0.4370 ;
        RECT 1.6470 0.0300 1.6970 0.4080 ;
        RECT 0.5830 0.0300 0.6330 0.5150 ;
        RECT 4.9910 0.0300 5.0410 0.2200 ;
        RECT 4.6870 0.0300 4.7370 0.3300 ;
        RECT 2.7570 0.0300 2.8070 0.2870 ;
        RECT 1.8020 0.1960 2.1530 0.2460 ;
        RECT 4.2150 0.3300 4.7530 0.3800 ;
        RECT 2.7570 0.2870 3.2170 0.3370 ;
        RECT 2.1030 0.2460 2.1530 0.4500 ;
        RECT 1.9510 0.2460 2.0010 0.4500 ;
        RECT 3.1670 0.3370 3.2170 0.4610 ;
        RECT 3.1670 0.2490 3.2170 0.2870 ;
        RECT 3.1670 0.1990 3.3920 0.2490 ;
    END
  END VSS

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2650 1.1610 5.3750 1.2210 ;
        RECT 5.1430 1.2210 5.3750 1.2710 ;
        RECT 5.3250 0.2040 5.3750 1.1610 ;
        RECT 5.1430 1.2710 5.1930 1.5460 ;
        RECT 5.1270 0.1540 5.3750 0.2040 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2360 1.3150 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 5.4720 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 4.9910 0.9470 5.0410 1.6420 ;
        RECT 4.7270 1.3580 4.7770 1.6420 ;
        RECT 3.3430 1.3280 3.3930 1.6420 ;
        RECT 1.6470 1.3640 1.6970 1.6420 ;
        RECT 4.0500 1.3080 4.7770 1.3580 ;
        RECT 3.1500 1.2780 3.3930 1.3280 ;
        RECT 1.6470 1.3140 2.1530 1.3640 ;
        RECT 1.9510 1.0980 2.0010 1.3140 ;
        RECT 2.1030 1.1110 2.1530 1.3140 ;
        RECT 1.6470 1.1340 1.6970 1.3140 ;
    END
  END VDD

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6800 0.7250 0.7300 ;
        RECT 0.4010 0.5530 0.5110 0.6800 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 0.6640 1.0110 0.8150 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9390 0.0880 4.0690 0.1380 ;
        RECT 3.9870 0.1380 4.0690 0.1640 ;
        RECT 2.9390 0.1380 3.0950 0.2070 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7690 1.4240 1.9410 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.1130 1.0090 5.2230 1.1190 ;
        RECT 5.1730 0.8540 5.2230 1.0090 ;
        RECT 4.8390 0.8040 5.2230 0.8540 ;
        RECT 4.8390 0.8540 4.8890 1.5460 ;
        RECT 5.1730 0.3590 5.2230 0.8040 ;
        RECT 4.8390 0.3090 5.2230 0.3590 ;
        RECT 4.8390 0.1480 4.8890 0.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q
  OBS
    LAYER PO ;
      RECT 2.4930 0.7900 2.5230 1.6060 ;
      RECT 4.6210 1.0120 4.6510 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 3.1010 0.0680 3.1310 0.6180 ;
      RECT 4.6210 0.0680 4.6510 0.7870 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 3.7090 0.8250 3.7390 1.6060 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 3.7090 0.0680 3.7390 0.6220 ;
      RECT 4.4690 0.0680 4.4990 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 3.1010 0.7580 3.1310 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 4.7730 0.0680 4.8030 1.6060 ;
      RECT 5.2290 0.0680 5.2590 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 4.3170 0.0680 4.3470 1.6060 ;
      RECT 5.0770 0.0680 5.1070 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 4.9250 0.0680 4.9550 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 2.4930 0.0680 2.5230 0.5420 ;
      RECT 5.3810 0.0680 5.4110 1.6060 ;
    LAYER NWELL ;
      RECT -0.1150 0.6790 5.5870 1.7730 ;
    LAYER M1 ;
      RECT 1.4520 0.6040 1.6370 0.6540 ;
      RECT 0.2050 0.8880 1.5020 0.9380 ;
      RECT 1.4520 0.6540 1.5020 0.8880 ;
      RECT 0.2050 0.5280 0.2550 0.8880 ;
      RECT 0.2050 0.4780 0.3290 0.5280 ;
      RECT 0.2790 0.3180 0.3290 0.4780 ;
      RECT 0.2790 0.9380 0.3290 1.2160 ;
      RECT 3.6230 0.5050 3.7130 0.5550 ;
      RECT 3.6630 0.5550 3.7130 1.0010 ;
      RECT 3.6230 0.4700 3.6730 0.5050 ;
      RECT 2.7660 1.0010 3.7130 1.0510 ;
      RECT 3.4400 0.4200 3.6730 0.4700 ;
      RECT 3.6230 1.0510 3.6730 1.3080 ;
      RECT 3.6230 0.3710 3.6730 0.4200 ;
      RECT 3.4710 1.3080 3.6730 1.3580 ;
      RECT 3.4710 1.1010 3.5210 1.3080 ;
      RECT 2.3010 0.0960 2.7070 0.1460 ;
      RECT 4.2710 0.6040 4.9810 0.6540 ;
      RECT 4.2710 0.6540 4.3210 0.9780 ;
      RECT 3.9100 0.9780 4.3210 1.0280 ;
      RECT 3.9100 0.5880 3.9600 0.9780 ;
      RECT 3.9100 0.5380 4.0170 0.5880 ;
      RECT 2.6350 1.4780 3.1570 1.5280 ;
      RECT 2.6350 1.5280 2.6850 1.5650 ;
      RECT 0.7350 1.0420 0.9370 1.0920 ;
      RECT 0.8870 1.0920 0.9370 1.2160 ;
      RECT 0.7350 1.0920 0.7850 1.2160 ;
      RECT 0.7190 0.5120 1.2570 0.5620 ;
      RECT 0.8870 0.3120 1.5450 0.3620 ;
      RECT 1.4950 0.3620 1.5450 0.3940 ;
      RECT 0.8870 0.3620 0.9370 0.3940 ;
      RECT 2.4830 1.4280 2.5330 1.5260 ;
      RECT 2.4830 1.3780 3.2930 1.4280 ;
      RECT 3.2430 1.4280 3.2930 1.5840 ;
      RECT 2.0010 1.5260 2.5330 1.5760 ;
      RECT 1.7990 0.6180 2.2450 0.6680 ;
      RECT 1.7990 0.6680 1.8490 0.9140 ;
      RECT 1.7990 0.4220 1.8490 0.6180 ;
      RECT 2.2550 0.5180 2.3810 0.5680 ;
      RECT 2.2550 0.3940 2.3050 0.5180 ;
      RECT 2.3310 0.5680 2.3810 0.7180 ;
      RECT 2.2550 0.7180 2.3810 0.7680 ;
      RECT 2.2550 0.7680 2.3050 0.9140 ;
      RECT 4.2900 1.4290 4.6770 1.4790 ;
      RECT 4.4540 0.7090 4.6770 0.7590 ;
      RECT 4.4540 0.7590 4.5040 1.0990 ;
      RECT 3.8990 1.0990 4.5040 1.1490 ;
      RECT 3.8990 1.1490 3.9490 1.2720 ;
      RECT 3.7230 1.2720 3.9490 1.3220 ;
      RECT 3.7230 1.3220 3.7730 1.5280 ;
      RECT 3.5310 1.5280 3.7730 1.5780 ;
      RECT 2.6950 1.2780 3.0810 1.3280 ;
      RECT 1.1750 1.0880 1.5610 1.1380 ;
      RECT 4.3070 0.0880 4.3570 0.2300 ;
      RECT 3.4650 0.2300 4.3570 0.2800 ;
      RECT 3.4650 0.2800 3.5150 0.3140 ;
      RECT 3.3140 0.3140 3.5150 0.3640 ;
      RECT 3.3140 0.3640 3.3640 0.5400 ;
      RECT 3.0750 0.5400 3.3640 0.5900 ;
      RECT 3.6830 0.1880 3.7650 0.2300 ;
      RECT 2.5590 0.6400 3.4610 0.6900 ;
      RECT 2.5590 0.6900 2.6090 1.1580 ;
      RECT 2.5590 0.4840 2.6090 0.6400 ;
      RECT 2.5590 1.2080 2.6090 1.3140 ;
      RECT 2.5590 0.3550 2.6090 0.4340 ;
      RECT 2.5590 1.1580 2.9290 1.2080 ;
      RECT 2.5590 0.4340 2.7770 0.4840 ;
      RECT 2.4070 0.2990 2.4970 0.3810 ;
      RECT 2.4310 0.3810 2.4810 0.9880 ;
      RECT 1.0230 0.9880 2.4810 1.0380 ;
      RECT 2.4070 1.0380 2.4570 1.3140 ;
      RECT 1.3430 0.4620 1.3930 0.5040 ;
      RECT 1.0230 0.4120 1.3930 0.4620 ;
      RECT 1.6500 0.7760 1.7000 0.9880 ;
      RECT 1.6500 0.7260 1.7370 0.7760 ;
      RECT 1.6870 0.5540 1.7370 0.7260 ;
      RECT 1.3430 0.5040 1.7370 0.5540 ;
      RECT 3.7750 0.4380 5.1170 0.4880 ;
      RECT 5.0670 0.4880 5.1170 0.7040 ;
      RECT 4.7270 0.7040 5.1170 0.7540 ;
      RECT 3.7750 0.4880 3.8250 1.1650 ;
      RECT 4.0780 0.4880 4.1280 0.7660 ;
      RECT 4.0780 0.7660 4.2210 0.8160 ;
      RECT 4.7270 0.7540 4.7770 1.2080 ;
      RECT 4.3670 1.2080 4.7770 1.2580 ;
      RECT 3.0750 0.7860 3.5970 0.8360 ;
      RECT 3.5470 0.6210 3.5970 0.7860 ;
  END
END SDFFNARX1_LVT

MACRO SDFFNARX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.776 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.5690 0.0970 5.6790 0.2070 ;
        RECT 5.6110 0.2070 5.6610 0.2700 ;
        RECT 5.2950 0.2700 5.6610 0.3200 ;
        RECT 5.2950 0.1480 5.3450 0.2700 ;
        RECT 5.6110 0.3200 5.6610 0.9180 ;
        RECT 5.2950 0.9180 5.6610 0.9680 ;
        RECT 5.2950 0.9680 5.3450 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 5.7760 0.0300 ;
        RECT 1.8020 0.0300 1.8520 0.1960 ;
        RECT 0.4310 0.0300 0.4810 0.4370 ;
        RECT 1.6470 0.0300 1.6970 0.4080 ;
        RECT 5.4470 0.0300 5.4970 0.2200 ;
        RECT 0.5830 0.0300 0.6330 0.5150 ;
        RECT 4.8390 0.0300 4.8890 0.4080 ;
        RECT 5.1430 0.0300 5.1930 0.3190 ;
        RECT 4.6870 0.0300 4.7370 0.3300 ;
        RECT 2.7570 0.0300 2.8070 0.2870 ;
        RECT 1.8020 0.1960 2.1530 0.2460 ;
        RECT 4.2150 0.3300 4.7530 0.3800 ;
        RECT 2.7570 0.2870 3.2170 0.3370 ;
        RECT 2.1030 0.2460 2.1530 0.4500 ;
        RECT 1.9510 0.2460 2.0010 0.4500 ;
        RECT 3.1670 0.3370 3.2170 0.4610 ;
        RECT 3.1670 0.2490 3.2170 0.2870 ;
        RECT 3.1670 0.1990 3.3920 0.2490 ;
    END
  END VSS

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2360 1.3150 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.9910 0.1480 5.0410 0.3940 ;
        RECT 4.9910 0.3940 5.5370 0.4440 ;
        RECT 5.4170 0.4440 5.5370 0.5110 ;
        RECT 5.4870 0.5110 5.5370 0.8040 ;
        RECT 4.9910 0.8040 5.5370 0.8540 ;
        RECT 4.9910 0.8540 5.0410 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 5.7760 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 4.8390 0.9120 4.8890 1.6420 ;
        RECT 5.1430 0.9600 5.1930 1.6420 ;
        RECT 5.4470 1.0520 5.4970 1.6420 ;
        RECT 4.7270 1.3580 4.7770 1.6420 ;
        RECT 3.3430 1.3280 3.3930 1.6420 ;
        RECT 1.6470 1.3640 1.6970 1.6420 ;
        RECT 4.0500 1.3080 4.7770 1.3580 ;
        RECT 3.1500 1.2780 3.3930 1.3280 ;
        RECT 1.6470 1.3140 2.1530 1.3640 ;
        RECT 1.9510 1.0980 2.0010 1.3140 ;
        RECT 2.1030 1.1110 2.1530 1.3140 ;
        RECT 1.6470 1.1340 1.6970 1.3140 ;
    END
  END VDD

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6800 0.7250 0.7300 ;
        RECT 0.4010 0.5530 0.5110 0.6800 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 0.6640 1.0110 0.8150 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9390 0.0880 4.0690 0.1380 ;
        RECT 3.9870 0.1380 4.0690 0.1740 ;
        RECT 2.9390 0.1380 3.0950 0.2070 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7690 1.4240 1.9410 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  OBS
    LAYER PO ;
      RECT 3.1010 0.7580 3.1310 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 4.7730 0.0680 4.8030 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 4.3170 0.0680 4.3470 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 5.3810 0.0680 5.4110 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 4.9250 0.0680 4.9550 1.6060 ;
      RECT 5.0770 0.0680 5.1070 1.6060 ;
      RECT 5.2290 0.0680 5.2590 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 2.4930 0.0680 2.5230 0.5420 ;
      RECT 2.4930 0.7900 2.5230 1.6060 ;
      RECT 4.6210 1.0120 4.6510 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 3.1010 0.0680 3.1310 0.6180 ;
      RECT 4.6210 0.0680 4.6510 0.7870 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 3.7090 0.8250 3.7390 1.6060 ;
      RECT 5.6850 0.0680 5.7150 1.6060 ;
      RECT 5.5330 0.0680 5.5630 1.6060 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 3.7090 0.0680 3.7390 0.6220 ;
      RECT 4.4690 0.0680 4.4990 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
    LAYER NWELL ;
      RECT -0.1150 0.6790 5.8910 1.7730 ;
    LAYER M1 ;
      RECT 5.2000 0.6040 5.4370 0.6540 ;
      RECT 4.0980 0.7660 4.2210 0.8160 ;
      RECT 4.0980 0.4880 4.1480 0.7660 ;
      RECT 3.7750 0.4380 4.4800 0.4880 ;
      RECT 4.4300 0.4880 4.4800 0.5030 ;
      RECT 3.7750 0.4880 3.8250 1.1650 ;
      RECT 4.7270 0.7540 4.7770 1.2080 ;
      RECT 4.3670 1.2080 4.7770 1.2580 ;
      RECT 4.4300 0.5030 5.2500 0.5530 ;
      RECT 5.2000 0.5530 5.2500 0.6040 ;
      RECT 5.2000 0.6540 5.2500 0.7040 ;
      RECT 4.7270 0.7040 5.2500 0.7540 ;
      RECT 3.0750 0.7860 3.5970 0.8360 ;
      RECT 3.5470 0.6210 3.5970 0.7860 ;
      RECT 1.4520 0.6040 1.6370 0.6540 ;
      RECT 0.2050 0.8880 1.5020 0.9380 ;
      RECT 1.4520 0.6540 1.5020 0.8880 ;
      RECT 0.2050 0.5280 0.2550 0.8880 ;
      RECT 0.2790 0.9380 0.3290 1.2160 ;
      RECT 0.2050 0.4780 0.3290 0.5280 ;
      RECT 0.2790 0.3180 0.3290 0.4780 ;
      RECT 3.6230 0.5050 3.7130 0.5550 ;
      RECT 3.6630 0.5550 3.7130 1.0010 ;
      RECT 3.6230 0.4700 3.6730 0.5050 ;
      RECT 2.7660 1.0010 3.7130 1.0510 ;
      RECT 3.4400 0.4200 3.6730 0.4700 ;
      RECT 3.6230 1.0510 3.6730 1.3080 ;
      RECT 3.6230 0.3710 3.6730 0.4200 ;
      RECT 3.4710 1.3080 3.6730 1.3580 ;
      RECT 3.4710 1.1010 3.5210 1.3080 ;
      RECT 2.3010 0.0960 2.7070 0.1460 ;
      RECT 4.2710 0.6040 5.1330 0.6540 ;
      RECT 4.2710 0.6540 4.3210 0.9780 ;
      RECT 3.9100 0.9780 4.3210 1.0280 ;
      RECT 3.9920 0.5880 4.0420 0.9780 ;
      RECT 3.9110 0.5380 4.0420 0.5880 ;
      RECT 2.6350 1.4780 3.1570 1.5280 ;
      RECT 2.6350 1.5280 2.6850 1.5650 ;
      RECT 0.7350 1.0420 0.9370 1.0920 ;
      RECT 0.8870 1.0920 0.9370 1.2160 ;
      RECT 0.7350 1.0920 0.7850 1.2160 ;
      RECT 0.7190 0.5120 1.2570 0.5620 ;
      RECT 0.8870 0.3120 1.5450 0.3620 ;
      RECT 1.4950 0.3620 1.5450 0.3940 ;
      RECT 0.8870 0.3620 0.9370 0.3940 ;
      RECT 2.4830 1.4280 2.5330 1.5260 ;
      RECT 2.4830 1.3780 3.2930 1.4280 ;
      RECT 3.2430 1.4280 3.2930 1.5840 ;
      RECT 2.0010 1.5260 2.5330 1.5760 ;
      RECT 1.7990 0.6180 2.2450 0.6680 ;
      RECT 1.7990 0.6680 1.8490 0.9140 ;
      RECT 1.7990 0.4220 1.8490 0.6180 ;
      RECT 2.2550 0.5180 2.3810 0.5680 ;
      RECT 2.2550 0.3940 2.3050 0.5180 ;
      RECT 2.3310 0.5680 2.3810 0.7180 ;
      RECT 2.2550 0.7180 2.3810 0.7680 ;
      RECT 2.2550 0.7680 2.3050 0.9140 ;
      RECT 4.2900 1.4290 4.6770 1.4790 ;
      RECT 4.4540 0.7090 4.6770 0.7590 ;
      RECT 4.4540 0.7590 4.5040 1.0990 ;
      RECT 3.8990 1.0990 4.5040 1.1490 ;
      RECT 3.8990 1.1490 3.9490 1.2720 ;
      RECT 3.7230 1.2720 3.9490 1.3220 ;
      RECT 3.7230 1.3220 3.7730 1.5280 ;
      RECT 3.5310 1.5280 3.7730 1.5780 ;
      RECT 2.6950 1.2780 3.0810 1.3280 ;
      RECT 1.1750 1.0880 1.5610 1.1380 ;
      RECT 4.3070 0.0880 4.3570 0.2300 ;
      RECT 3.4650 0.2300 4.3570 0.2800 ;
      RECT 3.6830 0.2800 3.7650 0.2900 ;
      RECT 3.4650 0.2800 3.5150 0.3140 ;
      RECT 3.3140 0.3140 3.5150 0.3640 ;
      RECT 3.3140 0.3640 3.3640 0.5400 ;
      RECT 3.0750 0.5400 3.3640 0.5900 ;
      RECT 3.6830 0.1880 3.7650 0.2300 ;
      RECT 2.5590 0.6400 3.4610 0.6900 ;
      RECT 2.5590 0.6900 2.6090 1.1580 ;
      RECT 2.5590 0.4840 2.6090 0.6400 ;
      RECT 2.5590 1.2080 2.6090 1.3140 ;
      RECT 2.5590 0.3550 2.6090 0.4340 ;
      RECT 2.5590 1.1580 2.9290 1.2080 ;
      RECT 2.5590 0.4340 2.7770 0.4840 ;
      RECT 2.4070 0.2990 2.4970 0.3810 ;
      RECT 2.4310 0.3810 2.4810 0.9880 ;
      RECT 1.0230 0.9880 2.4810 1.0380 ;
      RECT 2.4070 1.0380 2.4570 1.3140 ;
      RECT 1.3430 0.4620 1.3930 0.5040 ;
      RECT 1.0230 0.4120 1.3930 0.4620 ;
      RECT 1.6500 0.7760 1.7000 0.9880 ;
      RECT 1.6500 0.7260 1.7370 0.7760 ;
      RECT 1.6870 0.5540 1.7370 0.7260 ;
      RECT 1.3430 0.5040 1.7370 0.5540 ;
  END
END SDFFNARX2_LVT

MACRO SDFFNASRX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.776 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4170 1.0090 5.5270 1.1190 ;
        RECT 5.4770 0.8540 5.5270 1.0090 ;
        RECT 5.1430 0.8040 5.5270 0.8540 ;
        RECT 5.1430 0.8540 5.1930 1.5460 ;
        RECT 5.4770 0.3590 5.5270 0.8040 ;
        RECT 5.1430 0.3090 5.5270 0.3590 ;
        RECT 5.1430 0.1480 5.1930 0.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7690 1.4240 1.9410 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 5.7760 0.0300 ;
        RECT 1.6470 0.0300 1.6970 0.1960 ;
        RECT 0.5830 0.0300 0.6330 0.5150 ;
        RECT 5.2950 0.0300 5.3450 0.2200 ;
        RECT 0.4310 0.0300 0.4810 0.4370 ;
        RECT 2.7570 0.0300 2.8070 0.2870 ;
        RECT 4.9910 0.0300 5.0410 0.3300 ;
        RECT 1.6470 0.1960 2.1530 0.2460 ;
        RECT 2.7570 0.2870 3.3690 0.3370 ;
        RECT 4.3670 0.3300 5.0570 0.3800 ;
        RECT 1.9510 0.2460 2.0010 0.4500 ;
        RECT 2.1030 0.2460 2.1530 0.4500 ;
        RECT 1.6470 0.2460 1.6970 0.4080 ;
        RECT 3.1670 0.3370 3.2170 0.4610 ;
        RECT 3.3190 0.3370 3.3690 0.4610 ;
    END
  END VSS

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.7470 0.8570 4.9190 1.0340 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2360 1.3150 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6800 0.7250 0.7300 ;
        RECT 0.4010 0.5530 0.5110 0.6800 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9390 0.0880 4.2210 0.1380 ;
        RECT 4.1390 0.1380 4.2210 0.1640 ;
        RECT 2.9390 0.1380 3.0950 0.2070 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 0.6640 1.0110 0.8150 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 5.7760 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 5.2950 0.9470 5.3450 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 5.0310 1.3580 5.0810 1.6420 ;
        RECT 3.3430 1.3280 3.3930 1.6420 ;
        RECT 1.6470 1.3540 1.6970 1.6420 ;
        RECT 4.2020 1.3080 5.0810 1.3580 ;
        RECT 3.1500 1.2780 3.5520 1.3280 ;
        RECT 1.6470 1.3040 2.1530 1.3540 ;
        RECT 1.9510 1.0880 2.0010 1.3040 ;
        RECT 2.1030 1.0880 2.1530 1.3040 ;
        RECT 1.6470 1.1340 1.6970 1.3040 ;
    END
  END VDD

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.5690 1.1610 5.6790 1.2210 ;
        RECT 5.4470 1.2210 5.6790 1.2710 ;
        RECT 5.6290 0.2040 5.6790 1.1610 ;
        RECT 5.4470 1.2710 5.4970 1.5460 ;
        RECT 5.4310 0.1540 5.6790 0.2040 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN
  OBS
    LAYER PO ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 4.7730 0.0680 4.8030 1.6060 ;
      RECT 4.3170 0.0680 4.3470 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 5.5330 0.0680 5.5630 1.6060 ;
      RECT 5.0770 0.0680 5.1070 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 2.4930 0.0680 2.5230 0.4920 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 3.1010 0.8640 3.1310 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 4.9250 1.0120 4.9550 1.6060 ;
      RECT 3.8610 0.7320 3.8910 1.6060 ;
      RECT 3.8610 0.0680 3.8910 0.5820 ;
      RECT 3.1010 0.0680 3.1310 0.6680 ;
      RECT 4.9250 0.0680 4.9550 0.7870 ;
      RECT 2.4930 0.7900 2.5230 1.6060 ;
      RECT 5.6850 0.0680 5.7150 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 5.2290 0.0680 5.2590 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 4.6210 0.0680 4.6510 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 5.3810 0.0680 5.4110 1.6060 ;
      RECT 4.4690 0.0680 4.4990 1.6060 ;
      RECT 3.7090 0.0680 3.7390 1.6060 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
    LAYER NWELL ;
      RECT -0.1000 0.6790 5.9060 1.7730 ;
    LAYER M1 ;
      RECT 1.4520 0.6040 1.6370 0.6540 ;
      RECT 0.2050 0.5280 0.2550 0.8880 ;
      RECT 0.2790 0.9380 0.3290 1.2160 ;
      RECT 0.2050 0.4780 0.3290 0.5280 ;
      RECT 0.2790 0.3180 0.3290 0.4780 ;
      RECT 0.2050 0.8880 1.5020 0.9380 ;
      RECT 1.4520 0.6540 1.5020 0.8880 ;
      RECT 3.0750 0.8920 3.6640 0.9420 ;
      RECT 3.6140 0.7420 3.6640 0.8920 ;
      RECT 3.6140 0.6920 3.7650 0.7420 ;
      RECT 2.7660 1.0010 3.8650 1.0510 ;
      RECT 3.8150 0.6400 3.8650 1.0010 ;
      RECT 3.7750 1.0510 3.8250 1.3080 ;
      RECT 3.7750 0.5900 3.8650 0.6400 ;
      RECT 3.6230 1.3080 3.8250 1.3580 ;
      RECT 3.7750 0.4960 3.8250 0.5900 ;
      RECT 3.6230 1.2160 3.6730 1.3080 ;
      RECT 3.6230 0.4460 3.8250 0.4960 ;
      RECT 3.3020 1.1660 3.6730 1.2160 ;
      RECT 3.6230 0.3710 3.6730 0.4460 ;
      RECT 3.7750 0.3710 3.8250 0.4460 ;
      RECT 2.2550 0.4310 2.3810 0.4810 ;
      RECT 2.2550 0.1460 2.3050 0.4310 ;
      RECT 2.3310 0.4810 2.3810 0.8640 ;
      RECT 2.2550 0.0960 2.7070 0.1460 ;
      RECT 2.2320 0.8640 2.3810 0.9140 ;
      RECT 2.0030 1.5260 2.5330 1.5760 ;
      RECT 2.4830 1.4280 2.5330 1.5260 ;
      RECT 2.4830 1.3780 3.2930 1.4280 ;
      RECT 3.2430 1.4280 3.2930 1.5440 ;
      RECT 1.7990 0.5350 2.0770 0.5850 ;
      RECT 2.0270 0.5850 2.0770 0.7230 ;
      RECT 1.7990 0.5850 1.8490 0.9140 ;
      RECT 1.7990 0.4220 1.8490 0.5350 ;
      RECT 0.7350 1.0420 0.9370 1.0920 ;
      RECT 0.7350 1.0920 0.7850 1.2160 ;
      RECT 0.8870 1.0920 0.9370 1.2160 ;
      RECT 0.7190 0.5120 1.2570 0.5620 ;
      RECT 4.5610 0.7090 4.9810 0.7590 ;
      RECT 4.5610 0.7590 4.6110 1.0990 ;
      RECT 4.0510 1.0990 4.6110 1.1490 ;
      RECT 4.0510 1.1490 4.1010 1.2720 ;
      RECT 3.8750 1.2720 4.1010 1.3220 ;
      RECT 3.8750 1.3220 3.9250 1.4280 ;
      RECT 3.6830 1.4280 3.9250 1.4780 ;
      RECT 0.8870 0.3120 1.5450 0.3620 ;
      RECT 1.4950 0.3620 1.5450 0.3940 ;
      RECT 0.8870 0.3620 0.9370 0.3940 ;
      RECT 4.4230 0.6040 5.2850 0.6540 ;
      RECT 4.4230 0.6540 4.4730 0.9780 ;
      RECT 4.0620 0.9780 4.4730 1.0280 ;
      RECT 4.0620 0.5880 4.1120 0.9780 ;
      RECT 4.0620 0.5380 4.1690 0.5880 ;
      RECT 2.6350 1.4780 3.1570 1.5280 ;
      RECT 2.6350 1.5280 2.6850 1.5650 ;
      RECT 4.4420 1.4080 4.9810 1.4580 ;
      RECT 2.6950 1.2780 3.0810 1.3280 ;
      RECT 4.5190 1.2080 4.9050 1.2580 ;
      RECT 3.5020 1.5280 4.8420 1.5780 ;
      RECT 1.1750 1.0880 1.5610 1.1380 ;
      RECT 5.3710 0.4880 5.4210 0.7040 ;
      RECT 3.9270 0.4380 5.4210 0.4880 ;
      RECT 5.0310 0.7040 5.4210 0.7540 ;
      RECT 5.0310 0.7540 5.0810 1.1080 ;
      RECT 4.6710 1.1080 5.0810 1.1580 ;
      RECT 4.2300 0.4880 4.2800 0.7660 ;
      RECT 3.9270 0.4880 3.9770 1.1650 ;
      RECT 4.2300 0.7660 4.3730 0.8160 ;
      RECT 2.4070 0.2990 2.4970 0.3810 ;
      RECT 2.4310 0.3810 2.4810 0.9880 ;
      RECT 2.4070 1.0380 2.4570 1.3140 ;
      RECT 1.0230 0.9880 2.4810 1.0380 ;
      RECT 1.3430 0.4620 1.3930 0.5040 ;
      RECT 1.0230 0.4120 1.3930 0.4620 ;
      RECT 1.6500 0.7760 1.7000 0.9880 ;
      RECT 1.6500 0.7260 1.7370 0.7760 ;
      RECT 1.6870 0.5540 1.7370 0.7260 ;
      RECT 1.3430 0.5040 1.7370 0.5540 ;
      RECT 2.5590 0.7880 3.4610 0.8380 ;
      RECT 2.5590 0.4840 2.6090 0.7880 ;
      RECT 2.5590 0.8380 2.6090 1.1580 ;
      RECT 2.5590 0.3550 2.6090 0.4340 ;
      RECT 2.5590 1.2080 2.6090 1.3140 ;
      RECT 2.5590 0.4340 2.7770 0.4840 ;
      RECT 2.5590 1.1580 2.9290 1.2080 ;
      RECT 4.4590 0.0880 4.5090 0.2300 ;
      RECT 3.5110 0.2300 4.5090 0.2800 ;
      RECT 3.5110 0.2800 3.5610 0.5900 ;
      RECT 3.0750 0.5900 3.5610 0.6400 ;
      RECT 3.8350 0.1880 3.9170 0.2300 ;
  END
END SDFFNASRX1_LVT

MACRO SDFFNASRX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.08 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7690 1.4240 1.9410 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 6.0800 0.0300 ;
        RECT 1.6470 0.0300 1.6970 0.1960 ;
        RECT 0.4310 0.0300 0.4810 0.4370 ;
        RECT 5.1430 0.0300 5.1930 0.4080 ;
        RECT 0.5830 0.0300 0.6330 0.5150 ;
        RECT 5.7510 0.0300 5.8010 0.2200 ;
        RECT 5.4470 0.0300 5.4970 0.3190 ;
        RECT 2.7570 0.0300 2.8070 0.2870 ;
        RECT 4.9910 0.0300 5.0410 0.3300 ;
        RECT 1.6470 0.1960 2.1530 0.2460 ;
        RECT 2.7570 0.2870 3.3690 0.3370 ;
        RECT 4.3670 0.3300 5.0570 0.3800 ;
        RECT 1.9510 0.2460 2.0010 0.4500 ;
        RECT 2.1030 0.2460 2.1530 0.4500 ;
        RECT 1.6470 0.2460 1.6970 0.4080 ;
        RECT 3.1670 0.3370 3.2170 0.4610 ;
        RECT 3.3190 0.3370 3.3690 0.4610 ;
    END
  END VSS

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.7470 0.8570 4.9190 1.0340 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2360 1.3150 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6800 0.7250 0.7300 ;
        RECT 0.4010 0.5530 0.5110 0.6800 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9390 0.0880 4.2210 0.1380 ;
        RECT 4.1390 0.1380 4.2210 0.1740 ;
        RECT 2.9390 0.1380 3.0950 0.2070 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 0.6640 1.0110 0.8150 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 6.0800 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 5.4470 0.9600 5.4970 1.6420 ;
        RECT 5.1430 0.9120 5.1930 1.6420 ;
        RECT 5.7510 1.0520 5.8010 1.6420 ;
        RECT 5.0310 1.3580 5.0810 1.6420 ;
        RECT 3.3430 1.3280 3.3930 1.6420 ;
        RECT 1.6470 1.3540 1.6970 1.6420 ;
        RECT 4.2020 1.3080 5.0810 1.3580 ;
        RECT 3.1500 1.2780 3.5520 1.3280 ;
        RECT 1.6470 1.3040 2.1530 1.3540 ;
        RECT 1.9510 1.0880 2.0010 1.3040 ;
        RECT 2.1030 1.0880 2.1530 1.3040 ;
        RECT 1.6470 1.1340 1.6970 1.3040 ;
    END
  END VDD

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8730 0.0970 5.9830 0.2070 ;
        RECT 5.9150 0.2070 5.9650 0.2700 ;
        RECT 5.5990 0.2700 5.9650 0.3200 ;
        RECT 5.5990 0.1480 5.6490 0.2700 ;
        RECT 5.9150 0.3200 5.9650 0.9180 ;
        RECT 5.5990 0.9180 5.9650 0.9680 ;
        RECT 5.5990 0.9680 5.6490 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2950 0.8040 5.8410 0.8540 ;
        RECT 5.2950 0.8540 5.3450 1.5460 ;
        RECT 5.7910 0.5110 5.8410 0.8040 ;
        RECT 5.7210 0.4440 5.8410 0.5110 ;
        RECT 5.2950 0.3940 5.8410 0.4440 ;
        RECT 5.2950 0.1480 5.3450 0.3940 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q
  OBS
    LAYER PO ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 4.9250 1.0120 4.9550 1.6060 ;
      RECT 5.6850 0.0680 5.7150 1.6060 ;
      RECT 5.2290 0.0680 5.2590 1.6060 ;
      RECT 5.3810 0.0680 5.4110 1.6060 ;
      RECT 5.5330 0.0680 5.5630 1.6060 ;
      RECT 5.9890 0.0680 6.0190 1.6060 ;
      RECT 5.8370 0.0680 5.8670 1.6060 ;
      RECT 3.8610 0.7320 3.8910 1.6060 ;
      RECT 3.8610 0.0680 3.8910 0.5820 ;
      RECT 3.1010 0.0680 3.1310 0.6680 ;
      RECT 4.9250 0.0680 4.9550 0.7870 ;
      RECT 2.4930 0.7900 2.5230 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 4.6210 0.0680 4.6510 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 4.4690 0.0680 4.4990 1.6060 ;
      RECT 3.7090 0.0680 3.7390 1.6060 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 3.1010 0.8640 3.1310 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 4.7730 0.0680 4.8030 1.6060 ;
      RECT 4.3170 0.0680 4.3470 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 5.0770 0.0680 5.1070 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 2.4930 0.0680 2.5230 0.4920 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
    LAYER NWELL ;
      RECT -0.1000 0.6790 6.2100 1.7730 ;
    LAYER M1 ;
      RECT 2.5590 0.7880 3.4610 0.8380 ;
      RECT 2.5590 0.8380 2.6090 1.1580 ;
      RECT 2.5590 0.4840 2.6090 0.7880 ;
      RECT 2.5590 1.2080 2.6090 1.3140 ;
      RECT 2.5590 0.3550 2.6090 0.4340 ;
      RECT 2.5590 1.1580 2.9290 1.2080 ;
      RECT 2.5590 0.4340 2.7770 0.4840 ;
      RECT 4.4590 0.0880 4.5090 0.2300 ;
      RECT 3.5110 0.2300 4.5090 0.2800 ;
      RECT 3.8350 0.2800 3.9170 0.2900 ;
      RECT 3.5110 0.2800 3.5610 0.5900 ;
      RECT 3.0750 0.5900 3.5610 0.6400 ;
      RECT 3.8350 0.1880 3.9170 0.2300 ;
      RECT 1.4520 0.6040 1.6370 0.6540 ;
      RECT 0.2050 0.5280 0.2550 0.8880 ;
      RECT 0.2790 0.9380 0.3290 1.2160 ;
      RECT 0.2050 0.4780 0.3290 0.5280 ;
      RECT 0.2790 0.3180 0.3290 0.4780 ;
      RECT 0.2050 0.8880 1.5020 0.9380 ;
      RECT 1.4520 0.6540 1.5020 0.8880 ;
      RECT 3.0750 0.8920 3.6640 0.9420 ;
      RECT 3.6140 0.7420 3.6640 0.8920 ;
      RECT 3.6140 0.6920 3.7650 0.7420 ;
      RECT 3.7750 0.5900 3.8650 0.6400 ;
      RECT 3.8150 0.6400 3.8650 1.0010 ;
      RECT 3.7750 0.4960 3.8250 0.5900 ;
      RECT 2.7660 1.0010 3.8650 1.0510 ;
      RECT 3.6230 0.4460 3.8250 0.4960 ;
      RECT 3.7750 1.0510 3.8250 1.3080 ;
      RECT 3.6230 0.3710 3.6730 0.4460 ;
      RECT 3.7750 0.3710 3.8250 0.4460 ;
      RECT 3.6230 1.3080 3.8250 1.3580 ;
      RECT 3.6230 1.2160 3.6730 1.3080 ;
      RECT 3.3020 1.1660 3.6730 1.2160 ;
      RECT 2.2550 0.4310 2.3810 0.4810 ;
      RECT 2.2550 0.1460 2.3050 0.4310 ;
      RECT 2.3310 0.4810 2.3810 0.8640 ;
      RECT 2.2550 0.0960 2.7070 0.1460 ;
      RECT 2.2320 0.8640 2.3810 0.9140 ;
      RECT 2.0030 1.5260 2.5330 1.5760 ;
      RECT 2.4830 1.4280 2.5330 1.5260 ;
      RECT 2.4830 1.3780 3.2930 1.4280 ;
      RECT 3.2430 1.4280 3.2930 1.5440 ;
      RECT 1.7990 0.5350 2.0770 0.5850 ;
      RECT 2.0270 0.5850 2.0770 0.7230 ;
      RECT 1.7990 0.5850 1.8490 0.9140 ;
      RECT 1.7990 0.4220 1.8490 0.5350 ;
      RECT 0.7350 1.0420 0.9370 1.0920 ;
      RECT 0.7350 1.0920 0.7850 1.2160 ;
      RECT 0.8870 1.0920 0.9370 1.2160 ;
      RECT 0.7190 0.5120 1.2570 0.5620 ;
      RECT 4.5610 0.7090 4.9810 0.7590 ;
      RECT 4.5610 0.7590 4.6110 1.0990 ;
      RECT 4.0510 1.0990 4.6110 1.1490 ;
      RECT 4.0510 1.1490 4.1010 1.2720 ;
      RECT 3.8750 1.2720 4.1010 1.3220 ;
      RECT 3.8750 1.3220 3.9250 1.4280 ;
      RECT 3.6830 1.4280 3.9250 1.4780 ;
      RECT 0.8870 0.3120 1.5450 0.3620 ;
      RECT 1.4950 0.3620 1.5450 0.3940 ;
      RECT 0.8870 0.3620 0.9370 0.3940 ;
      RECT 4.4230 0.6040 5.4370 0.6540 ;
      RECT 4.4230 0.6540 4.4730 0.9780 ;
      RECT 4.0620 0.9780 4.4730 1.0280 ;
      RECT 4.0620 0.5880 4.1120 0.9780 ;
      RECT 4.0620 0.5380 4.1690 0.5880 ;
      RECT 2.6350 1.4780 3.1570 1.5280 ;
      RECT 2.6350 1.5280 2.6850 1.5650 ;
      RECT 4.4420 1.4080 4.9810 1.4580 ;
      RECT 2.6950 1.2780 3.0810 1.3280 ;
      RECT 4.5190 1.2080 4.9050 1.2580 ;
      RECT 3.5020 1.5280 4.8420 1.5780 ;
      RECT 1.1750 1.0880 1.5610 1.1380 ;
      RECT 5.5040 0.6040 5.7410 0.6540 ;
      RECT 5.0310 0.7540 5.0810 1.1080 ;
      RECT 4.6710 1.1080 5.0810 1.1580 ;
      RECT 4.5720 0.4880 4.6220 0.5030 ;
      RECT 3.9270 0.4380 4.6220 0.4880 ;
      RECT 3.9270 0.4880 3.9770 1.1650 ;
      RECT 4.2300 0.4880 4.2800 0.7660 ;
      RECT 4.2300 0.7660 4.3730 0.8160 ;
      RECT 5.5040 0.6540 5.5540 0.7040 ;
      RECT 5.5040 0.5530 5.5540 0.6040 ;
      RECT 4.5720 0.5030 5.5540 0.5530 ;
      RECT 5.0310 0.7040 5.5540 0.7540 ;
      RECT 2.4070 0.2990 2.4970 0.3810 ;
      RECT 2.4310 0.3810 2.4810 0.9880 ;
      RECT 2.4070 1.0380 2.4570 1.3140 ;
      RECT 1.0230 0.9880 2.4810 1.0380 ;
      RECT 1.3430 0.4620 1.3930 0.5040 ;
      RECT 1.0230 0.4120 1.3930 0.4620 ;
      RECT 1.6500 0.7760 1.7000 0.9880 ;
      RECT 1.6500 0.7260 1.7370 0.7760 ;
      RECT 1.6870 0.5540 1.7370 0.7260 ;
      RECT 1.3430 0.5040 1.7370 0.5540 ;
  END
END SDFFNASRX2_LVT

MACRO SDFFNASX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.472 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2360 1.3150 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6800 0.7250 0.7300 ;
        RECT 0.4010 0.5530 0.5110 0.6800 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2650 1.1610 5.3750 1.2210 ;
        RECT 5.1430 1.2210 5.3750 1.2710 ;
        RECT 5.3250 0.2040 5.3750 1.1610 ;
        RECT 5.1430 1.2710 5.1930 1.5460 ;
        RECT 5.1270 0.1540 5.3750 0.2040 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 0.6640 1.0110 0.8150 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 5.4720 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 4.9910 0.9470 5.0410 1.6420 ;
        RECT 3.1910 1.3210 3.2410 1.6420 ;
        RECT 4.7270 1.3580 4.7770 1.6420 ;
        RECT 1.6470 1.3600 1.6970 1.6420 ;
        RECT 2.9900 1.2710 3.4000 1.3210 ;
        RECT 4.0500 1.3080 4.7770 1.3580 ;
        RECT 1.6470 1.3100 2.1530 1.3600 ;
        RECT 1.9510 1.0940 2.0010 1.3100 ;
        RECT 2.1030 1.1070 2.1530 1.3100 ;
        RECT 1.6470 1.1340 1.6970 1.3100 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 5.4720 0.0300 ;
        RECT 1.8020 0.0300 1.8520 0.1960 ;
        RECT 0.4310 0.0300 0.4810 0.4370 ;
        RECT 0.5830 0.0300 0.6330 0.5150 ;
        RECT 3.1670 0.0300 3.2170 0.4610 ;
        RECT 4.9910 0.0300 5.0410 0.2200 ;
        RECT 1.6470 0.0300 1.6970 0.4080 ;
        RECT 3.0150 0.0300 3.0650 0.3710 ;
        RECT 4.6870 0.0300 4.7370 0.3300 ;
        RECT 1.8020 0.1960 2.1530 0.2460 ;
        RECT 4.0610 0.3300 4.7530 0.3800 ;
        RECT 2.1030 0.2460 2.1530 0.4500 ;
        RECT 1.9510 0.2460 2.0010 0.4500 ;
    END
  END VSS

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4430 0.8570 4.6150 1.0340 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7690 1.4240 1.9410 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.1130 1.0090 5.2230 1.1190 ;
        RECT 5.1730 0.8540 5.2230 1.0090 ;
        RECT 4.8390 0.8040 5.2230 0.8540 ;
        RECT 4.8390 0.8540 4.8890 1.5460 ;
        RECT 5.1730 0.3590 5.2230 0.8040 ;
        RECT 4.8390 0.3090 5.2230 0.3590 ;
        RECT 4.8390 0.1480 4.8890 0.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q
  OBS
    LAYER PO ;
      RECT 3.7090 0.7270 3.7390 1.6060 ;
      RECT 5.3810 0.0680 5.4110 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 2.4930 0.0680 2.5230 0.5420 ;
      RECT 3.1010 0.0660 3.1310 1.6040 ;
      RECT 4.6210 0.0680 4.6510 0.7870 ;
      RECT 4.0130 0.0650 4.0430 1.6030 ;
      RECT 2.7970 0.0660 2.8270 1.6040 ;
      RECT 2.6450 0.0660 2.6750 1.6040 ;
      RECT 2.9490 0.0660 2.9790 0.6620 ;
      RECT 2.4930 0.7900 2.5230 1.6060 ;
      RECT 4.6210 1.0120 4.6510 1.6060 ;
      RECT 2.9490 0.8300 2.9790 1.6040 ;
      RECT 3.7090 0.0680 3.7390 0.6220 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 4.7730 0.0680 4.8030 1.6060 ;
      RECT 5.2290 0.0680 5.2590 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 4.4690 0.0680 4.4990 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 5.0770 0.0680 5.1070 1.6060 ;
      RECT 4.3170 0.0680 4.3470 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 4.9250 0.0680 4.9550 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
    LAYER NWELL ;
      RECT -0.1150 0.6790 5.5870 1.7730 ;
    LAYER M1 ;
      RECT 2.7660 1.0010 3.7130 1.0510 ;
      RECT 3.6230 1.0510 3.6730 1.3080 ;
      RECT 3.6630 0.4960 3.7130 1.0010 ;
      RECT 3.4710 1.3080 3.6730 1.3580 ;
      RECT 3.4710 0.4460 3.7130 0.4960 ;
      RECT 3.4710 1.2160 3.5210 1.3080 ;
      RECT 3.6230 0.3710 3.6730 0.4460 ;
      RECT 3.4710 0.3710 3.5210 0.4460 ;
      RECT 3.1500 1.1660 3.5210 1.2160 ;
      RECT 4.2670 0.7090 4.6770 0.7590 ;
      RECT 4.2670 0.7590 4.3170 1.0990 ;
      RECT 3.8990 1.0990 4.3170 1.1490 ;
      RECT 3.8990 1.1490 3.9490 1.2720 ;
      RECT 3.8990 1.0960 3.9490 1.0990 ;
      RECT 3.7230 1.2720 3.9490 1.3220 ;
      RECT 3.7230 1.3220 3.7730 1.4280 ;
      RECT 3.5310 1.4280 3.7730 1.4780 ;
      RECT 0.7190 0.5120 1.2570 0.5620 ;
      RECT 0.8870 0.3120 1.5450 0.3620 ;
      RECT 1.4950 0.3620 1.5450 0.3940 ;
      RECT 0.8870 0.3620 0.9370 0.3940 ;
      RECT 4.1690 0.6040 4.9810 0.6050 ;
      RECT 4.1480 0.6050 4.9810 0.6540 ;
      RECT 4.1480 0.6540 4.1980 0.9750 ;
      RECT 3.8870 0.9750 4.1980 1.0240 ;
      RECT 3.8870 0.5850 3.9370 0.9750 ;
      RECT 3.9040 1.0240 4.1980 1.0250 ;
      RECT 3.8870 0.5350 3.9930 0.5850 ;
      RECT 2.6350 1.4760 3.0050 1.5260 ;
      RECT 2.6350 1.5260 2.6850 1.5630 ;
      RECT 2.0110 1.5260 2.5330 1.5760 ;
      RECT 2.4830 1.4260 2.5330 1.5260 ;
      RECT 2.4830 1.3760 3.1410 1.4260 ;
      RECT 3.0910 1.4260 3.1410 1.5410 ;
      RECT 4.1380 1.5190 4.6770 1.5690 ;
      RECT 1.7990 0.6180 2.2450 0.6680 ;
      RECT 1.7990 0.6680 1.8490 0.9140 ;
      RECT 1.7990 0.4220 1.8490 0.6180 ;
      RECT 2.2550 0.5180 2.3810 0.5680 ;
      RECT 2.2550 0.3940 2.3050 0.5180 ;
      RECT 2.3310 0.5680 2.3810 0.7180 ;
      RECT 2.2550 0.7180 2.3810 0.7680 ;
      RECT 2.2550 0.7680 2.3050 0.9140 ;
      RECT 3.3500 1.5280 3.8980 1.5780 ;
      RECT 3.8480 1.4610 3.8980 1.5280 ;
      RECT 3.8480 1.4110 4.5250 1.4610 ;
      RECT 2.3150 0.0960 2.7070 0.1460 ;
      RECT 0.7350 1.0420 0.9370 1.0920 ;
      RECT 0.8870 1.0920 0.9370 1.2160 ;
      RECT 0.7350 1.0920 0.7850 1.2160 ;
      RECT 1.1750 1.0880 1.5610 1.1380 ;
      RECT 4.2150 1.2080 4.6010 1.2580 ;
      RECT 4.1550 0.1490 4.2050 0.2300 ;
      RECT 3.3590 0.2300 4.2050 0.2800 ;
      RECT 3.6830 0.1780 3.7650 0.2300 ;
      RECT 3.3590 0.2800 3.4090 0.5840 ;
      RECT 2.9220 0.5840 3.4090 0.6340 ;
      RECT 3.3590 0.6340 3.4090 0.6360 ;
      RECT 2.4070 0.2990 2.4970 0.3810 ;
      RECT 2.4310 0.3810 2.4810 0.9880 ;
      RECT 1.0230 0.9880 2.4810 1.0380 ;
      RECT 2.4070 1.0380 2.4570 1.3140 ;
      RECT 1.3430 0.4620 1.3930 0.5040 ;
      RECT 1.0230 0.4120 1.3930 0.4620 ;
      RECT 1.6500 0.7760 1.7000 0.9880 ;
      RECT 1.6500 0.7260 1.7370 0.7760 ;
      RECT 1.6870 0.5540 1.7370 0.7260 ;
      RECT 1.3430 0.5040 1.7370 0.5540 ;
      RECT 5.0670 0.4810 5.1170 0.7040 ;
      RECT 3.7750 0.4310 5.1170 0.4810 ;
      RECT 4.7270 0.7040 5.1170 0.7540 ;
      RECT 4.7270 0.7540 4.7770 1.1080 ;
      RECT 4.3670 1.1080 4.7770 1.1580 ;
      RECT 3.7750 0.4810 3.8250 1.1650 ;
      RECT 4.0430 0.4810 4.0930 0.6960 ;
      RECT 3.9870 0.6960 4.0930 0.7460 ;
      RECT 2.9140 0.8780 3.5970 0.9280 ;
      RECT 3.5470 0.5970 3.5970 0.8780 ;
      RECT 1.4520 0.6040 1.6370 0.6540 ;
      RECT 0.2050 0.5280 0.2550 0.8880 ;
      RECT 0.2790 0.9380 0.3290 1.2160 ;
      RECT 0.2050 0.4780 0.3290 0.5280 ;
      RECT 0.2790 0.3180 0.3290 0.4780 ;
      RECT 0.2050 0.8880 1.5020 0.9380 ;
      RECT 1.4520 0.6540 1.5020 0.8880 ;
      RECT 2.5590 0.7440 3.3090 0.7940 ;
      RECT 2.5590 0.7940 2.6090 1.1560 ;
      RECT 2.5590 0.4820 2.6090 0.7440 ;
      RECT 2.5590 1.1560 2.7770 1.2060 ;
      RECT 2.5590 0.4320 2.7770 0.4820 ;
      RECT 2.5590 1.2060 2.6090 1.3140 ;
      RECT 2.5590 0.3550 2.6090 0.4320 ;
  END
END SDFFNASX1_LVT

MACRO SDFFNASX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.776 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2360 1.3150 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.5690 0.0970 5.6790 0.2070 ;
        RECT 5.6110 0.2070 5.6610 0.2700 ;
        RECT 5.2950 0.2700 5.6610 0.3200 ;
        RECT 5.2950 0.1480 5.3450 0.2700 ;
        RECT 5.6110 0.3200 5.6610 0.9180 ;
        RECT 5.2950 0.9180 5.6610 0.9680 ;
        RECT 5.2950 0.9680 5.3450 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6800 0.7250 0.7300 ;
        RECT 0.4010 0.5530 0.5110 0.6800 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.9910 0.8040 5.5370 0.8540 ;
        RECT 4.9910 0.8540 5.0410 1.5460 ;
        RECT 5.4870 0.5110 5.5370 0.8040 ;
        RECT 5.4170 0.4440 5.5370 0.5110 ;
        RECT 4.9910 0.3940 5.5370 0.4440 ;
        RECT 4.9910 0.1480 5.0410 0.3940 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 0.6640 1.0110 0.8150 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 5.7760 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 4.8390 0.9120 4.8890 1.6420 ;
        RECT 5.4470 1.0520 5.4970 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 5.1430 0.9600 5.1930 1.6420 ;
        RECT 4.7270 1.3580 4.7770 1.6420 ;
        RECT 3.1910 1.3210 3.2410 1.6420 ;
        RECT 1.6470 1.3600 1.6970 1.6420 ;
        RECT 4.0500 1.3080 4.7770 1.3580 ;
        RECT 2.9900 1.2710 3.4000 1.3210 ;
        RECT 1.6470 1.3100 2.1530 1.3600 ;
        RECT 1.9510 1.0940 2.0010 1.3100 ;
        RECT 2.1030 1.1070 2.1530 1.3100 ;
        RECT 1.6470 1.1340 1.6970 1.3100 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 5.7760 0.0300 ;
        RECT 1.8020 0.0300 1.8520 0.1960 ;
        RECT 0.4310 0.0300 0.4810 0.4370 ;
        RECT 0.5830 0.0300 0.6330 0.5150 ;
        RECT 4.8390 0.0300 4.8890 0.4080 ;
        RECT 5.4470 0.0300 5.4970 0.2200 ;
        RECT 5.1430 0.0300 5.1930 0.3190 ;
        RECT 3.1670 0.0300 3.2170 0.4610 ;
        RECT 1.6470 0.0300 1.6970 0.4080 ;
        RECT 3.0150 0.0300 3.0650 0.3710 ;
        RECT 4.6870 0.0300 4.7370 0.3300 ;
        RECT 1.8020 0.1960 2.1530 0.2460 ;
        RECT 4.0610 0.3300 4.7530 0.3800 ;
        RECT 2.1030 0.2460 2.1530 0.4500 ;
        RECT 1.9510 0.2460 2.0010 0.4500 ;
    END
  END VSS

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4430 0.8570 4.6150 1.0340 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7690 1.4240 1.9410 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  OBS
    LAYER PO ;
      RECT 2.4930 0.7900 2.5230 1.6060 ;
      RECT 5.5330 0.0680 5.5630 1.6060 ;
      RECT 5.3810 0.0680 5.4110 1.6060 ;
      RECT 5.6850 0.0680 5.7150 1.6060 ;
      RECT 5.2290 0.0680 5.2590 1.6060 ;
      RECT 5.0770 0.0680 5.1070 1.6060 ;
      RECT 4.9250 0.0680 4.9550 1.6060 ;
      RECT 4.6210 1.0120 4.6510 1.6060 ;
      RECT 2.9490 0.8300 2.9790 1.6040 ;
      RECT 3.7090 0.0680 3.7390 0.6220 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 4.7730 0.0680 4.8030 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 4.4690 0.0680 4.4990 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 4.3170 0.0680 4.3470 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 3.7090 0.7270 3.7390 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 2.4930 0.0680 2.5230 0.5420 ;
      RECT 3.1010 0.0660 3.1310 1.6040 ;
      RECT 4.6210 0.0680 4.6510 0.7870 ;
      RECT 4.0130 0.0650 4.0430 1.6030 ;
      RECT 2.7970 0.0660 2.8270 1.6040 ;
      RECT 2.6450 0.0660 2.6750 1.6040 ;
      RECT 2.9490 0.0660 2.9790 0.6620 ;
    LAYER NWELL ;
      RECT -0.1150 0.6790 5.8910 1.7730 ;
    LAYER M1 ;
      RECT 1.4520 0.6040 1.6370 0.6540 ;
      RECT 0.2050 0.5280 0.2550 0.8880 ;
      RECT 0.2790 0.9380 0.3290 1.2160 ;
      RECT 0.2050 0.4780 0.3290 0.5280 ;
      RECT 0.2790 0.3180 0.3290 0.4780 ;
      RECT 0.2050 0.8880 1.5020 0.9380 ;
      RECT 1.4520 0.6540 1.5020 0.8880 ;
      RECT 2.5590 0.7440 3.3090 0.7940 ;
      RECT 2.5590 0.7940 2.6090 1.1560 ;
      RECT 2.5590 0.4820 2.6090 0.7440 ;
      RECT 2.5590 1.1560 2.7770 1.2060 ;
      RECT 2.5590 0.4320 2.7770 0.4820 ;
      RECT 2.5590 1.2060 2.6090 1.3140 ;
      RECT 2.5590 0.3550 2.6090 0.4320 ;
      RECT 4.2670 0.7090 4.6770 0.7590 ;
      RECT 4.2670 0.7590 4.3170 1.0990 ;
      RECT 3.8990 1.0990 4.3170 1.1490 ;
      RECT 3.8990 1.0960 3.9490 1.0990 ;
      RECT 3.8990 1.1490 3.9490 1.2720 ;
      RECT 3.7230 1.2720 3.9490 1.3220 ;
      RECT 3.7230 1.3220 3.7730 1.4280 ;
      RECT 3.5310 1.4280 3.7730 1.4780 ;
      RECT 4.2150 1.2080 4.6010 1.2580 ;
      RECT 3.1500 1.1660 3.5210 1.2160 ;
      RECT 3.4710 1.2160 3.5210 1.3080 ;
      RECT 3.4710 1.3080 3.6730 1.3580 ;
      RECT 3.6230 1.0510 3.6730 1.3080 ;
      RECT 2.7660 1.0010 3.7130 1.0510 ;
      RECT 3.6630 0.4960 3.7130 1.0010 ;
      RECT 3.4710 0.4460 3.7130 0.4960 ;
      RECT 3.6230 0.3710 3.6730 0.4460 ;
      RECT 3.4710 0.3710 3.5210 0.4460 ;
      RECT 0.7190 0.5120 1.2570 0.5620 ;
      RECT 0.8870 0.3120 1.5450 0.3620 ;
      RECT 1.4950 0.3620 1.5450 0.3940 ;
      RECT 0.8870 0.3620 0.9370 0.3940 ;
      RECT 4.1690 0.6040 5.1340 0.6050 ;
      RECT 4.1480 0.6050 5.1340 0.6540 ;
      RECT 4.1480 0.6540 4.1980 0.9750 ;
      RECT 3.8870 0.9750 4.1980 1.0240 ;
      RECT 3.8870 0.5850 3.9370 0.9750 ;
      RECT 3.9040 1.0240 4.1980 1.0250 ;
      RECT 3.8870 0.5350 3.9930 0.5850 ;
      RECT 2.6350 1.4760 3.0050 1.5260 ;
      RECT 2.6350 1.5260 2.6850 1.5630 ;
      RECT 2.0110 1.5260 2.5330 1.5760 ;
      RECT 2.4830 1.4260 2.5330 1.5260 ;
      RECT 2.4830 1.3760 3.1410 1.4260 ;
      RECT 3.0910 1.4260 3.1410 1.5840 ;
      RECT 4.1380 1.5190 4.6770 1.5690 ;
      RECT 1.7990 0.6180 2.2450 0.6680 ;
      RECT 1.7990 0.6680 1.8490 0.9140 ;
      RECT 1.7990 0.4220 1.8490 0.6180 ;
      RECT 2.2550 0.5180 2.3810 0.5680 ;
      RECT 2.2550 0.3940 2.3050 0.5180 ;
      RECT 2.3310 0.5680 2.3810 0.7180 ;
      RECT 2.2550 0.7180 2.3810 0.7680 ;
      RECT 2.2550 0.7680 2.3050 0.9140 ;
      RECT 3.3500 1.5280 3.8980 1.5780 ;
      RECT 3.8480 1.4610 3.8980 1.5280 ;
      RECT 3.8480 1.4110 4.5250 1.4610 ;
      RECT 2.3150 0.0960 2.7070 0.1460 ;
      RECT 0.7350 1.0420 0.9370 1.0920 ;
      RECT 0.8870 1.0920 0.9370 1.2160 ;
      RECT 0.7350 1.0920 0.7850 1.2160 ;
      RECT 1.1750 1.0880 1.5610 1.1380 ;
      RECT 4.1550 0.0880 4.2050 0.2300 ;
      RECT 3.3590 0.2300 4.2050 0.2800 ;
      RECT 3.6830 0.1780 3.7650 0.2300 ;
      RECT 3.3590 0.2800 3.4090 0.5840 ;
      RECT 2.9220 0.5840 3.4090 0.6340 ;
      RECT 3.3590 0.6340 3.4090 0.6360 ;
      RECT 2.4070 0.2990 2.4970 0.3810 ;
      RECT 2.4310 0.3810 2.4810 0.9880 ;
      RECT 1.0230 0.9880 2.4810 1.0380 ;
      RECT 2.4070 1.0380 2.4570 1.3140 ;
      RECT 1.3430 0.4620 1.3930 0.5040 ;
      RECT 1.0230 0.4120 1.3930 0.4620 ;
      RECT 1.6500 0.7760 1.7000 0.9880 ;
      RECT 1.6500 0.7260 1.7370 0.7760 ;
      RECT 1.6870 0.5540 1.7370 0.7260 ;
      RECT 1.3430 0.5040 1.7370 0.5540 ;
      RECT 5.2000 0.6040 5.4370 0.6540 ;
      RECT 5.2000 0.5490 5.2500 0.6040 ;
      RECT 5.2000 0.6540 5.2500 0.7040 ;
      RECT 4.0430 0.4990 5.2500 0.5490 ;
      RECT 4.7270 0.7040 5.2500 0.7540 ;
      RECT 4.7270 0.7540 4.7770 1.1080 ;
      RECT 4.3670 1.1080 4.7770 1.1580 ;
      RECT 4.0430 0.5490 4.0930 0.6960 ;
      RECT 4.0430 0.4810 4.0930 0.4990 ;
      RECT 3.9870 0.6960 4.0930 0.7460 ;
      RECT 3.7750 0.4310 4.0930 0.4810 ;
      RECT 3.7750 0.4810 3.8250 1.1650 ;
      RECT 2.9140 0.8780 3.5970 0.9280 ;
      RECT 3.5470 0.5970 3.5970 0.8780 ;
  END
END SDFFNASX2_LVT

MACRO SDFFNX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.168 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.9610 1.1610 5.0710 1.2210 ;
        RECT 5.0210 0.2040 5.0710 1.1610 ;
        RECT 4.8390 1.2210 5.0710 1.2710 ;
        RECT 4.8230 0.1540 5.0710 0.2040 ;
        RECT 4.8390 1.2710 4.8890 1.5460 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8090 1.0090 4.9190 1.1190 ;
        RECT 4.8690 0.8540 4.9190 1.0090 ;
        RECT 4.5350 0.8040 4.9190 0.8540 ;
        RECT 4.5350 0.8540 4.5850 1.5460 ;
        RECT 4.8690 0.3590 4.9190 0.8040 ;
        RECT 4.5350 0.3090 4.9190 0.3590 ;
        RECT 4.5350 0.1480 4.5850 0.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7690 1.4240 1.9410 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 5.1680 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 4.6870 1.0190 4.7370 1.6420 ;
        RECT 4.4230 1.3580 4.4730 1.6420 ;
        RECT 3.8550 1.3580 3.9050 1.6420 ;
        RECT 3.1910 1.3280 3.2410 1.6420 ;
        RECT 1.6470 1.3540 1.6970 1.6420 ;
        RECT 4.3650 1.3080 4.4730 1.3580 ;
        RECT 3.8550 1.3080 3.9930 1.3580 ;
        RECT 2.9980 1.2780 3.2410 1.3280 ;
        RECT 1.6470 1.3040 2.1530 1.3540 ;
        RECT 2.1030 1.0880 2.1530 1.3040 ;
        RECT 1.9510 1.0880 2.0010 1.3040 ;
        RECT 1.6470 1.1340 1.6970 1.3040 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 0.6640 1.0110 0.8150 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6800 0.7250 0.7300 ;
        RECT 0.4010 0.5530 0.5110 0.6800 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2360 1.3150 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 5.1680 0.0300 ;
        RECT 1.6470 0.0300 1.6970 0.1960 ;
        RECT 3.0150 0.0300 3.0650 0.1990 ;
        RECT 4.6870 0.0300 4.7370 0.2200 ;
        RECT 0.5830 0.0300 0.6330 0.5150 ;
        RECT 0.4310 0.0300 0.4810 0.4370 ;
        RECT 4.3830 0.0300 4.4330 0.3300 ;
        RECT 1.6470 0.1960 2.1530 0.2460 ;
        RECT 3.0150 0.1990 3.2400 0.2490 ;
        RECT 3.9110 0.3300 4.4490 0.3800 ;
        RECT 2.1030 0.2460 2.1530 0.4500 ;
        RECT 1.9510 0.2460 2.0010 0.4500 ;
        RECT 1.6470 0.2460 1.6970 0.4080 ;
        RECT 3.0150 0.2490 3.0650 0.3730 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 5.2830 1.7730 ;
    LAYER M1 ;
      RECT 2.0110 1.5260 2.5330 1.5760 ;
      RECT 2.4830 1.4280 2.5330 1.5260 ;
      RECT 2.4830 1.3780 3.1410 1.4280 ;
      RECT 3.0910 1.4280 3.1410 1.5650 ;
      RECT 2.6350 1.4780 3.0050 1.5280 ;
      RECT 2.6350 1.5280 2.6850 1.5650 ;
      RECT 3.9860 1.5210 4.3730 1.5710 ;
      RECT 2.9230 0.7580 3.4450 0.8080 ;
      RECT 3.3950 0.5870 3.4450 0.7580 ;
      RECT 2.5590 0.6400 3.3090 0.6900 ;
      RECT 2.5590 0.4840 2.6090 0.6400 ;
      RECT 2.5590 0.6900 2.6090 1.1580 ;
      RECT 2.5590 0.4340 2.7770 0.4840 ;
      RECT 2.5590 1.1580 2.7770 1.2080 ;
      RECT 2.5590 0.3550 2.6090 0.4340 ;
      RECT 2.5590 1.2080 2.6090 1.3140 ;
      RECT 2.4070 0.2990 2.4970 0.3810 ;
      RECT 2.4310 0.3810 2.4810 0.9880 ;
      RECT 2.4070 1.0380 2.4570 1.3140 ;
      RECT 1.0230 0.9880 2.4810 1.0380 ;
      RECT 1.3430 0.4620 1.3930 0.5040 ;
      RECT 1.0230 0.4120 1.3930 0.4620 ;
      RECT 1.6500 0.7760 1.7000 0.9880 ;
      RECT 1.6500 0.7260 1.7370 0.7760 ;
      RECT 1.6870 0.5540 1.7370 0.7260 ;
      RECT 1.3430 0.5040 1.7370 0.5540 ;
      RECT 4.7630 0.4880 4.8130 0.7040 ;
      RECT 3.6230 0.4380 4.8130 0.4880 ;
      RECT 4.4230 0.7040 4.8130 0.7540 ;
      RECT 4.4230 0.7540 4.4730 1.2080 ;
      RECT 4.0630 1.2080 4.4730 1.2580 ;
      RECT 3.6230 0.4880 3.6730 1.1650 ;
      RECT 3.9260 0.4880 3.9760 0.6990 ;
      RECT 3.8350 0.6990 3.9760 0.7490 ;
      RECT 3.3310 0.1530 4.0530 0.2030 ;
      RECT 4.0030 0.2030 4.0530 0.2050 ;
      RECT 4.0030 0.1220 4.0530 0.1530 ;
      RECT 3.5310 0.1010 3.6130 0.1530 ;
      RECT 3.3310 0.2030 3.3810 0.3140 ;
      RECT 3.1800 0.3140 3.3810 0.3640 ;
      RECT 3.1800 0.3640 3.2300 0.5400 ;
      RECT 2.9230 0.5400 3.2300 0.5900 ;
      RECT 2.7660 1.0010 3.5610 1.0510 ;
      RECT 3.5110 0.4700 3.5610 1.0010 ;
      RECT 3.4710 1.0510 3.5210 1.3080 ;
      RECT 3.2880 0.4200 3.5610 0.4700 ;
      RECT 3.3190 1.3080 3.5210 1.3580 ;
      RECT 3.4710 0.3710 3.5210 0.4200 ;
      RECT 3.3190 1.1660 3.3690 1.3080 ;
      RECT 1.4520 0.6040 1.6370 0.6540 ;
      RECT 0.2050 0.5280 0.2550 0.8880 ;
      RECT 0.2790 0.9380 0.3290 1.2160 ;
      RECT 0.2050 0.4780 0.3290 0.5280 ;
      RECT 0.2790 0.3180 0.3290 0.4780 ;
      RECT 0.2050 0.8880 1.5020 0.9380 ;
      RECT 1.4520 0.6540 1.5020 0.8880 ;
      RECT 0.8870 0.3120 1.5450 0.3620 ;
      RECT 1.4950 0.3620 1.5450 0.3940 ;
      RECT 0.8870 0.3620 0.9370 0.3940 ;
      RECT 0.7190 0.5120 1.2570 0.5620 ;
      RECT 0.7350 1.0420 0.9370 1.0920 ;
      RECT 0.7350 1.0920 0.7850 1.2160 ;
      RECT 0.8870 1.0920 0.9370 1.2160 ;
      RECT 1.1750 1.0880 1.5610 1.1380 ;
      RECT 2.3150 0.0960 2.7070 0.1460 ;
      RECT 1.7990 0.6180 2.2450 0.6680 ;
      RECT 1.7990 0.6680 1.8490 0.9140 ;
      RECT 1.7990 0.4220 1.8490 0.6180 ;
      RECT 2.2550 0.5180 2.3810 0.5680 ;
      RECT 2.2550 0.3940 2.3050 0.5180 ;
      RECT 2.3310 0.5680 2.3810 0.7180 ;
      RECT 2.2550 0.7180 2.3810 0.7680 ;
      RECT 2.2550 0.7680 2.3050 0.9140 ;
      RECT 4.0400 0.6040 4.6770 0.6540 ;
      RECT 4.0400 0.6540 4.0900 0.9780 ;
      RECT 3.7350 0.9780 4.0900 1.0270 ;
      RECT 3.7350 0.5880 3.7850 0.9780 ;
      RECT 3.7580 1.0270 4.0900 1.0280 ;
      RECT 3.7350 0.5380 3.8650 0.5880 ;
      RECT 4.0400 1.0280 4.0900 1.0290 ;
      RECT 4.1500 0.7090 4.3730 0.7590 ;
      RECT 3.7470 1.1490 3.7970 1.2720 ;
      RECT 3.5710 1.2720 3.7970 1.3220 ;
      RECT 3.5710 1.3220 3.6210 1.5220 ;
      RECT 3.3790 1.5220 3.6210 1.5720 ;
      RECT 4.1500 0.7590 4.2000 1.0990 ;
      RECT 3.7470 1.0990 4.2000 1.1490 ;
    LAYER PO ;
      RECT 3.5570 0.7900 3.5870 1.6060 ;
      RECT 2.9490 0.0680 2.9790 0.6180 ;
      RECT 4.3170 0.0680 4.3470 0.7870 ;
      RECT 2.4930 0.7900 2.5230 1.6060 ;
      RECT 5.0770 0.0680 5.1070 1.6060 ;
      RECT 2.4930 0.0680 2.5230 0.5420 ;
      RECT 4.6210 0.0680 4.6510 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 4.7730 0.0680 4.8030 1.6060 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 3.7090 0.0680 3.7390 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 4.9250 0.0680 4.9550 1.6060 ;
      RECT 4.4690 0.0680 4.4990 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 2.9490 0.7300 2.9790 1.6060 ;
      RECT 3.5570 0.0680 3.5870 0.6220 ;
      RECT 4.3170 1.0120 4.3470 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
  END
END SDFFNX1_LVT

MACRO SDFFNX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.472 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2650 0.0970 5.3750 0.2070 ;
        RECT 5.3070 0.2070 5.3570 0.2700 ;
        RECT 4.9910 0.2700 5.3570 0.3200 ;
        RECT 4.9910 0.1480 5.0410 0.2700 ;
        RECT 5.3070 0.3200 5.3570 0.9180 ;
        RECT 4.9910 0.9180 5.3570 0.9680 ;
        RECT 4.9910 0.9680 5.0410 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7690 1.4240 1.9410 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 5.4720 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 4.8390 0.9600 4.8890 1.6420 ;
        RECT 4.5350 0.9120 4.5850 1.6420 ;
        RECT 5.1430 1.0520 5.1930 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 4.4230 1.3580 4.4730 1.6420 ;
        RECT 3.8550 1.3580 3.9050 1.6420 ;
        RECT 3.1910 1.3280 3.2410 1.6420 ;
        RECT 1.6470 1.3540 1.6970 1.6420 ;
        RECT 4.3650 1.3080 4.4730 1.3580 ;
        RECT 3.8550 1.3080 3.9930 1.3580 ;
        RECT 2.9980 1.2780 3.2410 1.3280 ;
        RECT 1.6470 1.3040 2.1530 1.3540 ;
        RECT 2.1030 1.0880 2.1530 1.3040 ;
        RECT 1.9510 1.0880 2.0010 1.3040 ;
        RECT 1.6470 1.1340 1.6970 1.3040 ;
    END
  END VDD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6870 0.1480 4.7370 0.3940 ;
        RECT 4.6870 0.3940 5.2330 0.4440 ;
        RECT 5.1130 0.4440 5.2330 0.5110 ;
        RECT 5.1830 0.5110 5.2330 0.8040 ;
        RECT 4.6870 0.8040 5.2330 0.8540 ;
        RECT 4.6870 0.8540 4.7370 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 0.6640 1.0110 0.8150 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6800 0.7250 0.7300 ;
        RECT 0.4010 0.5530 0.5110 0.6800 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2360 1.3150 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 5.4720 0.0300 ;
        RECT 1.6470 0.0300 1.6970 0.1960 ;
        RECT 3.0150 0.0300 3.0650 0.1990 ;
        RECT 0.4310 0.0300 0.4810 0.4370 ;
        RECT 4.5350 0.0300 4.5850 0.4080 ;
        RECT 5.1430 0.0300 5.1930 0.2200 ;
        RECT 4.8390 0.0300 4.8890 0.3190 ;
        RECT 0.5830 0.0300 0.6330 0.5150 ;
        RECT 4.3830 0.0300 4.4330 0.3300 ;
        RECT 1.6470 0.1960 2.1530 0.2460 ;
        RECT 3.0150 0.1990 3.2400 0.2490 ;
        RECT 3.9110 0.3300 4.4490 0.3800 ;
        RECT 2.1030 0.2460 2.1530 0.4500 ;
        RECT 1.9510 0.2460 2.0010 0.4500 ;
        RECT 1.6470 0.2460 1.6970 0.4080 ;
        RECT 3.0150 0.2490 3.0650 0.3730 ;
    END
  END VSS
  OBS
    LAYER PO ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 2.9490 0.7300 2.9790 1.6060 ;
      RECT 3.5570 0.0680 3.5870 0.6220 ;
      RECT 4.3170 1.0120 4.3470 1.6060 ;
      RECT 4.7730 0.0680 4.8030 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 4.6210 0.0680 4.6510 1.6060 ;
      RECT 3.5570 0.7900 3.5870 1.6060 ;
      RECT 2.9490 0.0680 2.9790 0.6180 ;
      RECT 4.3170 0.0680 4.3470 0.7870 ;
      RECT 2.4930 0.7900 2.5230 1.6060 ;
      RECT 5.3810 0.0680 5.4110 1.6060 ;
      RECT 2.4930 0.0680 2.5230 0.5420 ;
      RECT 5.2290 0.0680 5.2590 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 5.0770 0.0680 5.1070 1.6060 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 3.7090 0.0680 3.7390 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 4.9250 0.0680 4.9550 1.6060 ;
      RECT 4.4690 0.0680 4.4990 1.6060 ;
    LAYER NWELL ;
      RECT -0.1150 0.6790 5.5870 1.7730 ;
    LAYER M1 ;
      RECT 3.3310 0.1530 4.0530 0.2030 ;
      RECT 4.0030 0.0880 4.0530 0.1530 ;
      RECT 3.5310 0.1010 3.6130 0.1530 ;
      RECT 3.3310 0.2030 3.3810 0.3140 ;
      RECT 3.1800 0.3140 3.3810 0.3640 ;
      RECT 3.1800 0.3640 3.2300 0.5400 ;
      RECT 2.9230 0.5400 3.2300 0.5900 ;
      RECT 2.7660 1.0010 3.5610 1.0510 ;
      RECT 3.5110 0.4700 3.5610 1.0010 ;
      RECT 3.4710 1.0510 3.5210 1.3080 ;
      RECT 3.2880 0.4200 3.5610 0.4700 ;
      RECT 3.3190 1.3080 3.5210 1.3580 ;
      RECT 3.4710 0.3710 3.5210 0.4200 ;
      RECT 3.3190 1.1660 3.3690 1.3080 ;
      RECT 1.4520 0.6040 1.6370 0.6540 ;
      RECT 0.2050 0.5280 0.2550 0.8880 ;
      RECT 0.2790 0.9380 0.3290 1.2160 ;
      RECT 0.2050 0.4780 0.3290 0.5280 ;
      RECT 0.2790 0.3180 0.3290 0.4780 ;
      RECT 0.2050 0.8880 1.5020 0.9380 ;
      RECT 1.4520 0.6540 1.5020 0.8880 ;
      RECT 0.7350 1.0420 0.9370 1.0920 ;
      RECT 0.7350 1.0920 0.7850 1.2160 ;
      RECT 0.8870 1.0920 0.9370 1.2160 ;
      RECT 1.1750 1.0880 1.5610 1.1380 ;
      RECT 0.8870 0.3120 1.5450 0.3620 ;
      RECT 0.8870 0.3620 0.9370 0.3940 ;
      RECT 1.4950 0.3620 1.5450 0.3940 ;
      RECT 2.3150 0.0960 2.7070 0.1460 ;
      RECT 1.7990 0.6180 2.2450 0.6680 ;
      RECT 1.7990 0.6680 1.8490 0.9140 ;
      RECT 1.7990 0.4220 1.8490 0.6180 ;
      RECT 2.2550 0.5180 2.3810 0.5680 ;
      RECT 2.2550 0.3940 2.3050 0.5180 ;
      RECT 2.3310 0.5680 2.3810 0.7180 ;
      RECT 2.2550 0.7180 2.3810 0.7680 ;
      RECT 2.2550 0.7680 2.3050 0.9140 ;
      RECT 4.0400 0.6040 4.8290 0.6540 ;
      RECT 4.0400 0.6540 4.0900 0.9780 ;
      RECT 3.7350 0.9780 4.0900 1.0270 ;
      RECT 3.7350 0.5880 3.7850 0.9780 ;
      RECT 3.7580 1.0270 4.0900 1.0280 ;
      RECT 3.7350 0.5380 3.8650 0.5880 ;
      RECT 4.0400 1.0280 4.0900 1.0290 ;
      RECT 4.1500 0.7090 4.3730 0.7590 ;
      RECT 3.7470 1.1490 3.7970 1.2720 ;
      RECT 3.5710 1.2720 3.7970 1.3220 ;
      RECT 3.5710 1.3220 3.6210 1.5220 ;
      RECT 3.3790 1.5220 3.6210 1.5720 ;
      RECT 4.1500 0.7590 4.2000 1.0990 ;
      RECT 3.7470 1.0990 4.2000 1.1490 ;
      RECT 2.0110 1.5260 2.5330 1.5760 ;
      RECT 2.4830 1.4280 2.5330 1.5260 ;
      RECT 2.4830 1.3780 3.1410 1.4280 ;
      RECT 3.0910 1.4280 3.1410 1.5840 ;
      RECT 2.6350 1.4780 3.0050 1.5280 ;
      RECT 2.6350 1.5280 2.6850 1.5650 ;
      RECT 3.9860 1.5210 4.3730 1.5710 ;
      RECT 0.7190 0.5120 1.2570 0.5620 ;
      RECT 2.9230 0.7580 3.4450 0.8080 ;
      RECT 3.3950 0.5870 3.4450 0.7580 ;
      RECT 2.5590 0.6400 3.3090 0.6900 ;
      RECT 2.5590 0.4840 2.6090 0.6400 ;
      RECT 2.5590 0.6900 2.6090 1.1580 ;
      RECT 2.5590 0.4340 2.7770 0.4840 ;
      RECT 2.5590 1.1580 2.7770 1.2080 ;
      RECT 2.5590 0.3550 2.6090 0.4340 ;
      RECT 2.5590 1.2080 2.6090 1.3140 ;
      RECT 2.4070 0.2990 2.4970 0.3810 ;
      RECT 2.4310 0.3810 2.4810 0.9880 ;
      RECT 2.4070 1.0380 2.4570 1.3140 ;
      RECT 1.0230 0.9880 2.4810 1.0380 ;
      RECT 1.3430 0.4620 1.3930 0.5040 ;
      RECT 1.0230 0.4120 1.3930 0.4620 ;
      RECT 1.6500 0.7760 1.7000 0.9880 ;
      RECT 1.6500 0.7260 1.7370 0.7760 ;
      RECT 1.6870 0.5540 1.7370 0.7260 ;
      RECT 1.3430 0.5040 1.7370 0.5540 ;
      RECT 4.8960 0.6040 5.1330 0.6540 ;
      RECT 4.8960 0.5440 4.9460 0.6040 ;
      RECT 4.8960 0.6540 4.9460 0.7040 ;
      RECT 4.4230 0.7040 4.9460 0.7540 ;
      RECT 3.9260 0.4940 4.9460 0.5440 ;
      RECT 3.9260 0.5440 3.9760 0.6990 ;
      RECT 3.9260 0.4880 3.9760 0.4940 ;
      RECT 4.4230 0.7540 4.4730 1.2080 ;
      RECT 3.8350 0.6990 3.9760 0.7490 ;
      RECT 3.6230 0.4380 3.9760 0.4880 ;
      RECT 4.0630 1.2080 4.4730 1.2580 ;
      RECT 3.6230 0.4880 3.6730 1.1650 ;
  END
END SDFFNX2_LVT

MACRO RSDFFSRASRX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.336 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 10.3360 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 2.1030 1.1310 2.1530 1.6420 ;
        RECT 1.7990 1.1310 1.8490 1.6420 ;
        RECT 1.6470 1.1310 1.6970 1.6420 ;
        RECT 8.3750 1.4540 8.4250 1.6420 ;
        RECT 2.7110 1.2940 2.7610 1.6420 ;
        RECT 3.9670 1.2700 4.0170 1.6420 ;
        RECT 5.7510 1.4040 8.4250 1.4540 ;
        RECT 2.5390 1.2440 2.7610 1.2940 ;
        RECT 3.7580 1.2200 5.0570 1.2700 ;
        RECT 5.7510 1.2790 5.8010 1.4040 ;
        RECT 6.9670 0.9590 7.0170 1.4040 ;
        RECT 6.5110 0.9530 6.5610 1.4040 ;
    END
  END VDD

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.8150 0.4010 7.5150 0.4510 ;
        RECT 6.8150 0.1570 6.8650 0.4010 ;
        RECT 7.3930 0.4510 7.5150 0.5380 ;
        RECT 7.4650 0.5380 7.5150 0.8590 ;
        RECT 6.8150 0.8590 7.5150 0.9090 ;
        RECT 6.8150 0.9090 6.8650 1.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.1190 0.9690 7.6530 1.0190 ;
        RECT 7.6030 0.3510 7.6530 0.9690 ;
        RECT 7.1190 1.0190 7.3510 1.1290 ;
        RECT 7.1030 0.3010 7.6530 0.3510 ;
        RECT 7.1190 1.1290 7.1690 1.3270 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4670 1.4650 2.6390 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 10.3360 0.0300 ;
        RECT 2.1030 0.0300 2.1530 0.3070 ;
        RECT 9.3990 0.0300 9.4490 0.4260 ;
        RECT 1.6470 0.0300 1.6970 0.4050 ;
        RECT 6.9670 0.0300 7.0170 0.2410 ;
        RECT 1.7990 0.0300 1.8490 0.4050 ;
        RECT 8.0310 0.0300 8.0810 0.4260 ;
        RECT 0.5830 0.0300 0.6330 0.5120 ;
        RECT 0.4310 0.0300 0.4810 0.4340 ;
        RECT 8.9430 0.0300 8.9930 0.1980 ;
        RECT 6.6870 0.0300 6.7370 0.2930 ;
        RECT 2.1030 0.3070 3.9770 0.3570 ;
        RECT 5.7350 0.2930 6.7370 0.3400 ;
        RECT 2.5590 0.3570 2.6090 0.5570 ;
        RECT 3.7750 0.3570 3.8250 0.5570 ;
        RECT 2.7110 0.3570 2.7610 0.5570 ;
        RECT 3.9270 0.3570 3.9770 0.5330 ;
        RECT 2.1030 0.3570 2.1530 0.4050 ;
        RECT 3.9270 0.2440 3.9770 0.3070 ;
        RECT 5.7350 0.3400 6.7120 0.3430 ;
        RECT 3.9270 0.1940 5.0570 0.2440 ;
        RECT 4.3830 0.2440 4.4330 0.3490 ;
    END
  END VSS

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.9790 0.8570 6.1350 0.9750 ;
        RECT 5.9790 0.9750 6.0290 1.0790 ;
        RECT 5.4470 1.0790 6.0290 1.1290 ;
        RECT 5.4470 1.1290 5.4970 1.3200 ;
        RECT 4.1550 1.3200 5.4970 1.3700 ;
        RECT 4.1550 1.3700 4.2050 1.4550 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4390 0.0880 6.5120 0.1380 ;
        RECT 3.4390 0.1380 3.5970 0.2100 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.5210 0.2490 9.6310 0.3590 ;
        RECT 9.5320 0.3590 9.5820 0.5270 ;
        RECT 9.3070 0.5270 9.5820 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6570 0.7050 4.8130 0.7310 ;
        RECT 4.6570 0.7310 5.1170 0.7810 ;
        RECT 4.7630 0.5970 4.8130 0.7050 ;
        RECT 4.6570 0.7810 4.8130 0.8150 ;
        RECT 5.0670 0.7810 5.1170 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 8.0150 0.9470 9.6330 1.0070 ;
        RECT 9.5230 0.6900 9.6330 0.9470 ;
        RECT 9.3990 0.6270 9.4490 0.9470 ;
    END
  END VDDG

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2520 1.3330 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6780 0.7250 0.7280 ;
        RECT 0.4010 0.5510 0.5110 0.6780 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 1.1610 1.0110 1.3160 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D
  OBS
    LAYER M1 ;
      RECT 5.2950 1.0170 5.3450 1.1200 ;
      RECT 5.2950 1.1700 5.3450 1.2700 ;
      RECT 4.8230 1.1200 5.3450 1.1700 ;
      RECT 4.2130 0.8580 4.3730 0.9080 ;
      RECT 4.2130 0.9080 4.2630 0.9680 ;
      RECT 3.6830 0.9680 4.2630 1.0180 ;
      RECT 1.4520 0.6020 1.6370 0.6520 ;
      RECT 0.2050 0.8410 1.5020 0.8910 ;
      RECT 1.4520 0.6520 1.5020 0.8410 ;
      RECT 0.2050 0.5260 0.2550 0.8410 ;
      RECT 0.2790 0.8910 0.3290 1.2140 ;
      RECT 0.2050 0.4760 0.3290 0.5260 ;
      RECT 0.2790 0.3160 0.3290 0.4760 ;
      RECT 3.1670 0.8540 4.0690 0.9040 ;
      RECT 3.1670 0.6130 3.2170 0.8540 ;
      RECT 3.1670 0.9040 3.2170 1.0590 ;
      RECT 3.1670 0.5630 3.3690 0.6130 ;
      RECT 3.1670 1.0590 3.5370 1.1090 ;
      RECT 3.3190 0.4070 3.3690 0.5630 ;
      RECT 3.1670 0.4130 3.2170 0.5630 ;
      RECT 3.1670 1.1090 3.2170 1.3370 ;
      RECT 6.5870 0.6320 6.9410 0.6820 ;
      RECT 6.8910 0.5970 6.9410 0.6320 ;
      RECT 6.2590 0.7790 6.3090 1.1790 ;
      RECT 5.9430 0.7290 6.3090 0.7790 ;
      RECT 5.9430 0.4500 5.9930 0.7290 ;
      RECT 5.5990 0.4000 6.6370 0.4500 ;
      RECT 6.5870 0.4500 6.6370 0.6320 ;
      RECT 5.6000 1.1790 6.3090 1.2290 ;
      RECT 5.6000 1.2290 5.6500 1.3530 ;
      RECT 5.5990 0.4500 5.6490 0.5630 ;
      RECT 5.5990 0.2970 5.6490 0.4000 ;
      RECT 6.9910 0.6130 7.4130 0.6630 ;
      RECT 6.3590 0.8090 6.4090 1.3010 ;
      RECT 6.3590 0.5500 6.4090 0.7590 ;
      RECT 6.1310 0.5000 6.4090 0.5500 ;
      RECT 6.1310 0.5500 6.1810 0.6790 ;
      RECT 6.6630 0.8090 6.7130 1.3010 ;
      RECT 6.9910 0.6630 7.0410 0.7590 ;
      RECT 6.3590 0.7590 7.0410 0.8090 ;
      RECT 5.1470 0.1880 5.7410 0.2380 ;
      RECT 5.1470 0.2380 5.1970 0.2940 ;
      RECT 4.5060 0.2940 5.1970 0.3440 ;
      RECT 4.1190 0.4550 4.1690 0.6130 ;
      RECT 3.6830 0.6130 4.1690 0.6630 ;
      RECT 4.5060 0.3440 4.5560 0.4050 ;
      RECT 4.1190 0.4050 4.5560 0.4550 ;
      RECT 3.0150 0.8130 3.1050 0.8630 ;
      RECT 3.0550 0.4620 3.1050 0.8130 ;
      RECT 3.0150 0.8630 3.0650 1.0830 ;
      RECT 2.9990 0.4120 3.1050 0.4620 ;
      RECT 2.2550 1.0830 3.0650 1.1330 ;
      RECT 3.0150 1.1330 3.0650 1.3540 ;
      RECT 2.2550 0.7520 2.3050 1.0830 ;
      RECT 2.2550 0.7020 2.3450 0.7520 ;
      RECT 2.2950 0.5510 2.3450 0.7020 ;
      RECT 2.2550 0.5010 2.3450 0.5510 ;
      RECT 2.2550 0.4070 2.3050 0.5010 ;
      RECT 2.4070 0.6130 2.8530 0.6630 ;
      RECT 2.4070 0.6630 2.4570 1.0040 ;
      RECT 2.4070 0.4130 2.4570 0.6130 ;
      RECT 2.6180 0.0940 3.3150 0.1440 ;
      RECT 8.3190 0.8200 8.8670 0.8700 ;
      RECT 1.6500 0.7020 1.9410 0.7280 ;
      RECT 1.6870 0.6780 1.9410 0.7020 ;
      RECT 1.3430 0.4600 1.3930 0.5020 ;
      RECT 1.0230 0.4100 1.3930 0.4600 ;
      RECT 1.0230 1.0200 1.7000 1.0700 ;
      RECT 1.6500 0.7520 1.7000 1.0200 ;
      RECT 1.6500 0.7280 1.7370 0.7520 ;
      RECT 1.6870 0.5520 1.7370 0.6780 ;
      RECT 1.3430 0.5020 1.7370 0.5520 ;
      RECT 0.8870 0.3100 1.5450 0.3600 ;
      RECT 1.4950 0.3600 1.5450 0.3920 ;
      RECT 0.8870 0.3600 0.9370 0.3920 ;
      RECT 5.6590 0.8660 5.8080 0.9160 ;
      RECT 5.7580 0.9160 5.8080 0.9670 ;
      RECT 5.7580 0.9670 5.8930 1.0170 ;
      RECT 1.9910 0.6280 2.2450 0.6520 ;
      RECT 1.9520 0.6020 2.2450 0.6280 ;
      RECT 1.9910 0.6520 2.0410 0.7780 ;
      RECT 1.9520 0.5780 2.0410 0.6020 ;
      RECT 1.9520 0.7780 2.0410 0.8280 ;
      RECT 1.9520 0.3190 2.0020 0.5780 ;
      RECT 1.9520 0.8280 2.0020 1.0760 ;
      RECT 8.6230 0.7090 9.1610 0.7590 ;
      RECT 5.2010 1.5200 8.3250 1.5700 ;
      RECT 5.1830 0.5440 5.2330 1.0200 ;
      RECT 4.6710 0.5170 5.2330 0.5440 ;
      RECT 4.6870 1.0200 5.2330 1.0700 ;
      RECT 4.6710 0.4940 5.2320 0.5170 ;
      RECT 4.4230 0.7880 4.4730 1.1200 ;
      RECT 3.3740 0.7380 4.4750 0.7880 ;
      RECT 4.2310 0.5050 4.2810 0.7380 ;
      RECT 4.6870 1.0700 4.7370 1.1200 ;
      RECT 3.9110 1.1200 4.7370 1.1700 ;
      RECT 9.2470 0.6770 9.2970 0.7680 ;
      RECT 9.2070 0.4270 9.2970 0.4620 ;
      RECT 9.2470 0.1260 9.2970 0.4270 ;
      RECT 9.2070 0.6270 9.2970 0.6770 ;
      RECT 9.2070 0.5120 9.2570 0.6270 ;
      RECT 9.0030 0.4770 9.2570 0.5120 ;
      RECT 9.0030 0.4620 9.2970 0.4770 ;
      RECT 4.4430 1.5200 5.1330 1.5700 ;
      RECT 4.8980 0.6130 5.1330 0.6630 ;
      RECT 5.4470 0.8670 5.5890 0.9170 ;
      RECT 5.4470 0.6630 5.4970 0.8670 ;
      RECT 5.4470 0.6130 5.8930 0.6630 ;
      RECT 4.5350 0.9200 4.9650 0.9700 ;
      RECT 4.9150 0.8310 4.9650 0.9200 ;
      RECT 4.5350 0.9700 4.5850 1.0340 ;
      RECT 4.5350 0.5050 4.5850 0.9200 ;
      RECT 4.2910 1.4200 5.5970 1.4700 ;
      RECT 3.3030 1.1900 3.6890 1.2400 ;
      RECT 5.8800 1.2870 6.2730 1.3370 ;
      RECT 3.2270 1.3890 3.7650 1.4390 ;
      RECT 7.3310 1.2580 8.6290 1.3080 ;
      RECT 7.9390 0.5270 8.5370 0.5770 ;
      RECT 8.4870 0.5770 8.5370 0.7700 ;
      RECT 8.4870 0.3480 8.5370 0.5270 ;
      RECT 8.1830 0.5770 8.2330 0.8870 ;
      RECT 8.1830 0.1260 8.2330 0.5270 ;
      RECT 8.6230 0.1320 8.8570 0.1820 ;
      RECT 7.8790 1.1160 8.3280 1.1660 ;
      RECT 7.8790 0.6770 7.9290 1.1160 ;
      RECT 7.8390 0.6270 7.9290 0.6770 ;
      RECT 7.8390 0.4770 7.8890 0.6270 ;
      RECT 7.8390 0.4270 7.9290 0.4770 ;
      RECT 7.8790 0.1260 7.9290 0.4270 ;
      RECT 2.9230 1.5240 3.9170 1.5740 ;
      RECT 0.7190 0.5100 1.2570 0.5600 ;
      RECT 1.1750 1.1330 1.5610 1.1830 ;
      RECT 0.7190 0.9410 0.9530 0.9910 ;
      RECT 8.8510 1.1160 9.3890 1.1660 ;
      RECT 8.3190 0.2480 9.1610 0.2980 ;
      RECT 2.8630 0.7130 2.9890 0.7630 ;
      RECT 2.8630 0.7630 2.9130 1.0330 ;
      RECT 2.9390 0.5630 2.9890 0.7130 ;
      RECT 2.8470 0.5130 2.9890 0.5630 ;
      RECT 4.8230 0.3940 5.4970 0.4440 ;
      RECT 5.4470 0.4440 5.4970 0.5630 ;
      RECT 5.4470 0.2970 5.4970 0.3940 ;
      RECT 5.2950 0.9670 5.5130 1.0170 ;
      RECT 5.2950 0.4440 5.3450 0.9670 ;
    LAYER PO ;
      RECT 5.0770 0.8390 5.1070 1.6060 ;
      RECT 9.4850 0.0660 9.5150 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 5.8370 0.0660 5.8670 0.6910 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 3.1010 0.8400 3.1310 1.6060 ;
      RECT 5.8370 0.9390 5.8670 1.6060 ;
      RECT 5.5330 0.0660 5.5630 0.6370 ;
      RECT 3.1010 0.0660 3.1310 0.6370 ;
      RECT 9.3330 0.0660 9.3630 1.6060 ;
      RECT 3.7090 0.0660 3.7390 0.6910 ;
      RECT 5.0770 0.0660 5.1070 0.6910 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 9.6370 0.0660 9.6670 1.6060 ;
      RECT 4.7730 0.8920 4.8030 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 5.5330 0.8390 5.5630 1.6060 ;
      RECT 9.7890 0.0660 9.8190 1.6060 ;
      RECT 10.2450 0.0660 10.2750 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 9.9410 0.0660 9.9710 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 10.0930 0.0660 10.1230 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 4.7730 0.0660 4.8030 0.6910 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 3.7090 0.9390 3.7390 1.6060 ;
      RECT 7.3570 0.0670 7.3870 1.6050 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
    LAYER NWELL ;
      RECT 7.7120 0.4910 9.7230 1.0830 ;
      RECT -0.1150 1.5430 10.4580 1.7730 ;
      RECT -0.1150 0.6790 7.2500 1.5430 ;
      RECT 10.1830 0.6790 10.4580 1.5430 ;
  END
END RSDFFSRASRX1_LVT

MACRO RSDFFSRASRX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.64 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 10.6400 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 1.6470 1.1310 1.6970 1.6420 ;
        RECT 2.1030 1.1310 2.1530 1.6420 ;
        RECT 1.7990 1.1310 1.8490 1.6420 ;
        RECT 2.7110 1.2940 2.7610 1.6420 ;
        RECT 3.9670 1.2700 4.0170 1.6420 ;
        RECT 8.6790 1.4540 8.7290 1.6420 ;
        RECT 2.5390 1.2440 2.7610 1.2940 ;
        RECT 3.7580 1.2200 5.0570 1.2700 ;
        RECT 5.7510 1.4040 8.7290 1.4540 ;
        RECT 5.7510 1.2790 5.8010 1.4040 ;
        RECT 6.8150 0.9130 6.8650 1.4040 ;
        RECT 7.1190 0.9610 7.1690 1.4040 ;
        RECT 6.5110 0.9530 6.5610 1.4040 ;
        RECT 7.4230 1.0530 7.4730 1.4040 ;
    END
  END VDD

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4670 1.4650 2.6390 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0280 10.6400 0.0320 ;
        RECT 2.1030 0.0320 2.1530 0.3070 ;
        RECT 1.6470 0.0320 1.6970 0.4050 ;
        RECT 0.5830 0.0320 0.6330 0.5120 ;
        RECT 0.4310 0.0320 0.4810 0.4340 ;
        RECT 1.7990 0.0320 1.8490 0.4050 ;
        RECT 6.8150 0.0320 6.8650 0.4090 ;
        RECT 7.1190 0.0320 7.1690 0.3200 ;
        RECT 7.4230 0.0320 7.4730 0.2210 ;
        RECT 8.3350 0.0320 8.3850 0.4260 ;
        RECT 9.7030 0.0320 9.7530 0.4260 ;
        RECT 9.2470 0.0320 9.2970 0.1980 ;
        RECT 6.6870 0.0320 6.7370 0.2880 ;
        RECT 2.1030 0.3070 3.9770 0.3570 ;
        RECT 5.7350 0.2880 6.7370 0.3380 ;
        RECT 3.7750 0.3570 3.8250 0.5570 ;
        RECT 2.5590 0.3570 2.6090 0.5570 ;
        RECT 2.7110 0.3570 2.7610 0.5570 ;
        RECT 3.9270 0.3570 3.9770 0.5330 ;
        RECT 2.1030 0.3570 2.1530 0.4050 ;
        RECT 3.9270 0.2380 3.9770 0.3070 ;
        RECT 3.9270 0.1880 5.0570 0.2380 ;
        RECT 4.3830 0.2380 4.4330 0.3490 ;
    END
  END VSS

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.9790 0.8570 6.1350 0.9750 ;
        RECT 5.9790 0.9750 6.0290 1.0790 ;
        RECT 5.4470 1.0790 6.0290 1.1290 ;
        RECT 5.4470 1.1290 5.4970 1.3200 ;
        RECT 4.1550 1.3200 5.4970 1.3700 ;
        RECT 4.1550 1.3700 4.2050 1.4550 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END SETB

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.5470 0.0880 6.4850 0.0970 ;
        RECT 3.4390 0.0970 6.4850 0.1380 ;
        RECT 3.4390 0.1380 3.5970 0.2100 ;
        RECT 6.4350 0.1380 6.4850 0.1700 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.8250 0.2490 9.9350 0.3590 ;
        RECT 9.8360 0.3590 9.8860 0.5270 ;
        RECT 9.6110 0.5270 9.8860 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.7630 0.5970 4.8130 0.7050 ;
        RECT 4.6570 0.7050 4.8130 0.7310 ;
        RECT 4.6570 0.7310 5.1170 0.7810 ;
        RECT 4.6570 0.7810 4.8130 0.8150 ;
        RECT 5.0670 0.7810 5.1170 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.2710 0.1490 7.3210 0.2710 ;
        RECT 7.2710 0.2710 7.9690 0.3210 ;
        RECT 7.8460 0.3210 7.9690 0.3600 ;
        RECT 7.8460 0.2500 7.9690 0.2710 ;
        RECT 7.9190 0.3600 7.9690 0.9420 ;
        RECT 7.8460 0.2490 7.9610 0.2500 ;
        RECT 7.2710 0.9420 7.9690 0.9920 ;
        RECT 7.2710 0.9920 7.3210 1.3270 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 8.3190 0.9470 9.9370 1.0070 ;
        RECT 9.8270 0.6900 9.9370 0.9470 ;
        RECT 9.7030 0.6270 9.7530 0.9470 ;
    END
  END VDDG

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2520 1.3330 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6780 0.7250 0.7280 ;
        RECT 0.4010 0.5510 0.5110 0.6780 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.9670 0.8420 7.8190 0.8920 ;
        RECT 6.9670 0.8920 7.0170 1.3190 ;
        RECT 7.7690 0.5120 7.8190 0.8420 ;
        RECT 7.6970 0.4520 7.8190 0.5120 ;
        RECT 6.9670 0.4020 7.8190 0.4520 ;
        RECT 6.9670 0.1490 7.0170 0.4020 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 1.1610 1.0110 1.3160 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D
  OBS
    LAYER M1 ;
      RECT 5.2010 1.5200 8.6290 1.5700 ;
      RECT 1.4520 0.6020 1.6370 0.6520 ;
      RECT 0.2050 0.8410 1.5020 0.8910 ;
      RECT 1.4520 0.6520 1.5020 0.8410 ;
      RECT 0.2050 0.5260 0.2550 0.8410 ;
      RECT 0.2790 0.8910 0.3290 1.2140 ;
      RECT 0.2050 0.4760 0.3290 0.5260 ;
      RECT 0.2790 0.3160 0.3290 0.4760 ;
      RECT 0.8870 0.3100 1.5450 0.3600 ;
      RECT 1.4950 0.3600 1.5450 0.3920 ;
      RECT 0.8870 0.3600 0.9370 0.3920 ;
      RECT 1.6870 0.6780 1.9410 0.7020 ;
      RECT 1.6500 0.7020 1.9410 0.7280 ;
      RECT 1.3430 0.4600 1.3930 0.5020 ;
      RECT 1.0230 0.4100 1.3930 0.4600 ;
      RECT 1.3430 0.5020 1.7370 0.5520 ;
      RECT 1.6870 0.5520 1.7370 0.6780 ;
      RECT 1.6500 0.7280 1.7370 0.7520 ;
      RECT 1.6500 0.7520 1.7000 1.0200 ;
      RECT 1.0230 1.0200 1.7000 1.0700 ;
      RECT 0.7190 0.5100 1.2570 0.5600 ;
      RECT 3.1670 0.8540 4.0690 0.9040 ;
      RECT 3.1670 0.6130 3.2170 0.8540 ;
      RECT 3.1670 0.5630 3.3690 0.6130 ;
      RECT 3.1670 0.9040 3.2170 1.0590 ;
      RECT 3.3190 0.4070 3.3690 0.5630 ;
      RECT 3.1670 0.4130 3.2170 0.5630 ;
      RECT 3.1670 1.0590 3.5370 1.1090 ;
      RECT 3.1670 1.1090 3.2170 1.3370 ;
      RECT 1.9910 0.6280 2.2450 0.6520 ;
      RECT 1.9520 0.6020 2.2450 0.6280 ;
      RECT 1.9910 0.6520 2.0410 0.7780 ;
      RECT 1.9520 0.5780 2.0410 0.6020 ;
      RECT 1.9520 0.7780 2.0410 0.8280 ;
      RECT 1.9520 0.3190 2.0020 0.5780 ;
      RECT 1.9520 0.8280 2.0020 1.0760 ;
      RECT 2.8470 0.5130 2.9890 0.5630 ;
      RECT 2.9390 0.5630 2.9890 0.7130 ;
      RECT 2.8630 0.7130 2.9890 0.7630 ;
      RECT 2.8630 0.7630 2.9130 1.0330 ;
      RECT 2.9990 0.4120 3.1050 0.4620 ;
      RECT 3.0550 0.4620 3.1050 0.8130 ;
      RECT 3.0150 0.8130 3.1050 0.8630 ;
      RECT 3.0150 0.8630 3.0650 1.0830 ;
      RECT 2.2550 1.0830 3.0650 1.1330 ;
      RECT 3.0150 1.1330 3.0650 1.3540 ;
      RECT 2.2550 0.7520 2.3050 1.0830 ;
      RECT 2.2550 0.7020 2.3450 0.7520 ;
      RECT 2.2950 0.5510 2.3450 0.7020 ;
      RECT 2.2550 0.5010 2.3450 0.5510 ;
      RECT 2.2550 0.4070 2.3050 0.5010 ;
      RECT 2.4070 0.6130 2.8530 0.6630 ;
      RECT 2.4070 0.6630 2.4570 1.0040 ;
      RECT 2.4070 0.4130 2.4570 0.6130 ;
      RECT 2.6180 0.0940 3.3150 0.1440 ;
      RECT 5.1470 0.1880 5.7410 0.2380 ;
      RECT 5.1470 0.2380 5.1970 0.2880 ;
      RECT 4.5060 0.2880 5.1970 0.3380 ;
      RECT 4.1190 0.4550 4.1690 0.6130 ;
      RECT 3.6830 0.6130 4.1690 0.6630 ;
      RECT 4.5060 0.3380 4.5560 0.4050 ;
      RECT 4.1190 0.4050 4.5560 0.4550 ;
      RECT 4.8230 0.3880 5.4970 0.4380 ;
      RECT 5.4470 0.4380 5.4970 0.5630 ;
      RECT 5.4470 0.2970 5.4970 0.3880 ;
      RECT 5.2950 0.9670 5.5130 1.0170 ;
      RECT 5.2950 0.3840 5.3450 0.3880 ;
      RECT 5.2950 0.4380 5.3450 0.9670 ;
      RECT 5.2950 1.0170 5.3450 1.1200 ;
      RECT 5.2950 1.1700 5.3450 1.2700 ;
      RECT 4.8230 1.1200 5.3450 1.1700 ;
      RECT 6.5870 0.6420 7.1090 0.6920 ;
      RECT 5.9430 0.4500 5.9930 0.7290 ;
      RECT 5.9430 0.7290 6.3090 0.7790 ;
      RECT 6.2590 0.7790 6.3090 1.1790 ;
      RECT 6.5870 0.4500 6.6370 0.6420 ;
      RECT 5.5990 0.4000 6.6370 0.4500 ;
      RECT 5.6000 1.1790 6.3090 1.2290 ;
      RECT 5.5990 0.4500 5.6490 0.5630 ;
      RECT 5.5990 0.2970 5.6490 0.4000 ;
      RECT 5.6000 1.2290 5.6500 1.3530 ;
      RECT 4.6710 0.4880 5.2330 0.5380 ;
      RECT 5.1830 0.5380 5.2330 1.0200 ;
      RECT 4.6870 1.0200 5.2330 1.0700 ;
      RECT 4.4230 0.7880 4.4730 1.1200 ;
      RECT 3.3740 0.7380 4.4750 0.7880 ;
      RECT 4.2310 0.5050 4.2810 0.7380 ;
      RECT 4.6870 1.0700 4.7370 1.1200 ;
      RECT 3.9110 1.1200 4.7370 1.1700 ;
      RECT 4.8980 0.6130 5.1330 0.6630 ;
      RECT 5.4470 0.6130 5.8930 0.6630 ;
      RECT 5.4470 0.6630 5.4970 0.8670 ;
      RECT 5.4470 0.8670 5.5890 0.9170 ;
      RECT 4.5350 0.9200 4.9650 0.9700 ;
      RECT 4.9150 0.8310 4.9650 0.9200 ;
      RECT 4.5350 0.9700 4.5850 1.0340 ;
      RECT 4.5350 0.5050 4.5850 0.9200 ;
      RECT 7.1730 0.6130 7.7170 0.6630 ;
      RECT 6.3590 0.7920 6.4090 1.3010 ;
      RECT 6.3590 0.5500 6.4090 0.7420 ;
      RECT 6.1310 0.5000 6.4090 0.5500 ;
      RECT 6.1310 0.5500 6.1810 0.6790 ;
      RECT 6.6630 0.7920 6.7130 1.3010 ;
      RECT 7.1730 0.6630 7.2230 0.7420 ;
      RECT 6.3590 0.7420 7.2230 0.7920 ;
      RECT 8.1850 1.1070 8.6340 1.1170 ;
      RECT 8.1830 1.0670 8.6340 1.1070 ;
      RECT 8.1830 0.6770 8.2330 1.0670 ;
      RECT 8.1430 0.6270 8.2330 0.6770 ;
      RECT 8.1430 0.4770 8.1930 0.6270 ;
      RECT 8.1430 0.4270 8.2330 0.4770 ;
      RECT 8.1830 0.1260 8.2330 0.4270 ;
      RECT 8.2430 0.5270 8.8410 0.5770 ;
      RECT 8.7910 0.5770 8.8410 0.7700 ;
      RECT 8.7910 0.3480 8.8410 0.5270 ;
      RECT 8.4870 0.5770 8.5370 0.8870 ;
      RECT 8.4870 0.1260 8.5370 0.5270 ;
      RECT 8.6230 0.2480 9.4650 0.2980 ;
      RECT 9.5510 0.6770 9.6010 0.7680 ;
      RECT 9.5110 0.4270 9.6010 0.4620 ;
      RECT 9.5510 0.1260 9.6010 0.4270 ;
      RECT 9.5110 0.6270 9.6010 0.6770 ;
      RECT 9.5110 0.5120 9.5610 0.6270 ;
      RECT 9.3070 0.4770 9.5610 0.5120 ;
      RECT 9.3070 0.4620 9.6010 0.4770 ;
      RECT 8.9270 0.1320 9.1610 0.1820 ;
      RECT 1.1750 1.1330 1.5610 1.1830 ;
      RECT 0.7190 0.9410 0.9530 0.9910 ;
      RECT 3.3030 1.1900 3.6890 1.2400 ;
      RECT 3.2270 1.3890 3.7650 1.4390 ;
      RECT 3.6830 0.9680 4.2630 1.0180 ;
      RECT 4.2130 0.9080 4.2630 0.9680 ;
      RECT 4.2130 0.8580 4.3730 0.9080 ;
      RECT 2.9230 1.5240 3.9170 1.5740 ;
      RECT 5.7580 0.9670 5.8930 1.0170 ;
      RECT 5.7580 0.9160 5.8080 0.9670 ;
      RECT 5.6590 0.8660 5.8080 0.9160 ;
      RECT 4.4430 1.5200 5.1330 1.5700 ;
      RECT 4.2910 1.4200 5.5970 1.4700 ;
      RECT 5.8800 1.2870 6.2730 1.3370 ;
      RECT 7.6350 1.1990 8.9330 1.2490 ;
      RECT 8.6230 0.8200 9.1710 0.8700 ;
      RECT 8.9270 0.7090 9.4650 0.7590 ;
      RECT 9.1550 1.0670 9.6940 1.1170 ;
    LAYER PO ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 4.7730 0.0660 4.8030 0.6910 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 3.7090 0.9390 3.7390 1.6060 ;
      RECT 7.6610 0.0670 7.6910 1.6050 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 9.3330 0.0660 9.3630 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 5.0770 0.8390 5.1070 1.6060 ;
      RECT 9.7890 0.0660 9.8190 1.6060 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 9.4850 0.0660 9.5150 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 5.8370 0.0660 5.8670 0.6910 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 3.1010 0.8400 3.1310 1.6060 ;
      RECT 5.8370 0.9390 5.8670 1.6060 ;
      RECT 5.5330 0.0660 5.5630 0.6370 ;
      RECT 3.7090 0.0660 3.7390 0.6910 ;
      RECT 3.1010 0.0660 3.1310 0.6370 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 9.6370 0.0660 9.6670 1.6060 ;
      RECT 5.0770 0.0660 5.1070 0.6910 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 9.9410 0.0660 9.9710 1.6060 ;
      RECT 4.7730 0.8920 4.8030 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 5.5330 0.8390 5.5630 1.6060 ;
      RECT 10.0930 0.0660 10.1230 1.6060 ;
      RECT 10.5490 0.0660 10.5790 1.6060 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 10.2450 0.0660 10.2750 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 10.3970 0.0660 10.4270 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
    LAYER NWELL ;
      RECT 8.0160 0.4910 10.0270 1.0830 ;
      RECT -0.1150 1.5430 10.7620 1.7730 ;
      RECT -0.1150 0.6790 7.5540 1.5430 ;
      RECT 10.4870 0.6790 10.7620 1.5430 ;
  END
END RSDFFSRASRX2_LVT

MACRO RSDFFSRASX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.336 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 10.3360 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 2.1030 1.1310 2.1530 1.6420 ;
        RECT 1.7990 1.1310 1.8490 1.6420 ;
        RECT 1.6470 1.1310 1.6970 1.6420 ;
        RECT 8.3750 1.4540 8.4250 1.6420 ;
        RECT 2.7110 1.2940 2.7610 1.6420 ;
        RECT 3.9670 1.2700 4.0170 1.6420 ;
        RECT 5.7510 1.4040 8.4250 1.4540 ;
        RECT 2.5390 1.2440 2.7610 1.2940 ;
        RECT 3.7580 1.2200 5.0570 1.2700 ;
        RECT 5.7510 1.2790 5.8010 1.4040 ;
        RECT 6.9670 0.9590 7.0170 1.4040 ;
        RECT 6.5110 0.9530 6.5610 1.4040 ;
    END
  END VDD

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.8150 0.4010 7.5150 0.4510 ;
        RECT 6.8150 0.1570 6.8650 0.4010 ;
        RECT 7.3930 0.4510 7.5150 0.5380 ;
        RECT 7.4650 0.5380 7.5150 0.8590 ;
        RECT 6.8150 0.8590 7.5150 0.9090 ;
        RECT 6.8150 0.9090 6.8650 1.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.1190 0.9690 7.6530 1.0190 ;
        RECT 7.6030 0.3510 7.6530 0.9690 ;
        RECT 7.1190 1.0190 7.3510 1.1290 ;
        RECT 7.1030 0.3010 7.6530 0.3510 ;
        RECT 7.1190 1.1290 7.1690 1.3270 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4670 1.4650 2.6390 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 10.3360 0.0300 ;
        RECT 2.1030 0.0300 2.1530 0.3070 ;
        RECT 9.3990 0.0300 9.4490 0.4260 ;
        RECT 1.6470 0.0300 1.6970 0.4050 ;
        RECT 6.9670 0.0300 7.0170 0.2410 ;
        RECT 1.7990 0.0300 1.8490 0.4050 ;
        RECT 8.0310 0.0300 8.0810 0.4260 ;
        RECT 0.5830 0.0300 0.6330 0.5120 ;
        RECT 0.4310 0.0300 0.4810 0.4340 ;
        RECT 8.9430 0.0300 8.9930 0.1980 ;
        RECT 6.6870 0.0300 6.7370 0.2880 ;
        RECT 2.1030 0.3070 3.9770 0.3570 ;
        RECT 5.7350 0.2880 6.7370 0.3380 ;
        RECT 2.5590 0.3570 2.6090 0.5570 ;
        RECT 3.7750 0.3570 3.8250 0.5570 ;
        RECT 2.7110 0.3570 2.7610 0.5570 ;
        RECT 3.9270 0.3570 3.9770 0.5330 ;
        RECT 2.1030 0.3570 2.1530 0.4050 ;
        RECT 3.9270 0.2380 3.9770 0.3070 ;
        RECT 3.9270 0.1880 5.0570 0.2380 ;
        RECT 4.3830 0.2380 4.4330 0.3490 ;
    END
  END VSS

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.9790 0.8570 6.1350 0.9750 ;
        RECT 5.9790 0.9750 6.0290 1.0790 ;
        RECT 5.4470 1.0790 6.0290 1.1290 ;
        RECT 5.4470 1.1290 5.4970 1.3200 ;
        RECT 4.1550 1.3200 5.4970 1.3700 ;
        RECT 4.1550 1.3700 4.2050 1.4550 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.5210 0.2490 9.6310 0.3590 ;
        RECT 9.5320 0.3590 9.5820 0.5270 ;
        RECT 9.3070 0.5270 9.5820 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6570 0.7050 4.8130 0.7310 ;
        RECT 4.6570 0.7310 5.1170 0.7810 ;
        RECT 4.7630 0.5970 4.8130 0.7050 ;
        RECT 4.6570 0.7810 4.8130 0.8150 ;
        RECT 5.0670 0.7810 5.1170 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 8.0150 0.9470 9.6330 1.0070 ;
        RECT 9.5230 0.6900 9.6330 0.9470 ;
        RECT 9.3990 0.6270 9.4490 0.9470 ;
    END
  END VDDG

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2520 1.3330 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6780 0.7250 0.7280 ;
        RECT 0.4010 0.5510 0.5110 0.6780 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 1.1610 1.0110 1.3160 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D
  OBS
    LAYER M1 ;
      RECT 5.2950 0.9670 5.5130 1.0170 ;
      RECT 5.2950 0.4380 5.3450 0.9670 ;
      RECT 5.2950 1.0170 5.3450 1.1200 ;
      RECT 5.2950 1.1700 5.3450 1.2700 ;
      RECT 4.8230 1.1200 5.3450 1.1700 ;
      RECT 4.2130 0.8580 4.3730 0.9080 ;
      RECT 4.2130 0.9080 4.2630 0.9680 ;
      RECT 3.6830 0.9680 4.2630 1.0180 ;
      RECT 1.4520 0.6020 1.6370 0.6520 ;
      RECT 0.2050 0.8410 1.5020 0.8910 ;
      RECT 1.4520 0.6520 1.5020 0.8410 ;
      RECT 0.2050 0.5260 0.2550 0.8410 ;
      RECT 0.2790 0.8910 0.3290 1.2140 ;
      RECT 0.2050 0.4760 0.3290 0.5260 ;
      RECT 0.2790 0.3160 0.3290 0.4760 ;
      RECT 3.1670 0.8540 4.0690 0.9040 ;
      RECT 3.1670 0.6130 3.2170 0.8540 ;
      RECT 3.1670 0.9040 3.2170 1.0590 ;
      RECT 3.1670 0.5630 3.3690 0.6130 ;
      RECT 3.1670 1.0590 3.5370 1.1090 ;
      RECT 3.3190 0.4070 3.3690 0.5630 ;
      RECT 3.1670 0.4130 3.2170 0.5630 ;
      RECT 3.1670 1.1090 3.2170 1.3370 ;
      RECT 6.5600 0.6320 6.9410 0.6820 ;
      RECT 6.8910 0.5970 6.9410 0.6320 ;
      RECT 5.9430 0.4500 5.9930 0.7290 ;
      RECT 5.9430 0.7290 6.3090 0.7790 ;
      RECT 6.2590 0.7790 6.3090 1.1790 ;
      RECT 5.5990 0.4000 6.6370 0.4500 ;
      RECT 6.5870 0.4500 6.6370 0.6320 ;
      RECT 5.6000 1.1790 6.3090 1.2290 ;
      RECT 5.5990 0.4500 5.6490 0.5630 ;
      RECT 5.5990 0.2970 5.6490 0.4000 ;
      RECT 5.6000 1.2290 5.6500 1.3530 ;
      RECT 6.9910 0.6130 7.4130 0.6630 ;
      RECT 6.3590 0.8090 6.4090 1.3010 ;
      RECT 6.3590 0.5500 6.4090 0.7590 ;
      RECT 6.1310 0.5000 6.4090 0.5500 ;
      RECT 6.1310 0.5500 6.1810 0.6790 ;
      RECT 6.6630 0.8090 6.7130 1.3010 ;
      RECT 6.9910 0.6630 7.0410 0.7590 ;
      RECT 6.3590 0.7590 7.0410 0.8090 ;
      RECT 5.1470 0.1880 5.7410 0.2380 ;
      RECT 5.1470 0.2380 5.1970 0.2880 ;
      RECT 4.5060 0.2880 5.1970 0.3380 ;
      RECT 4.1190 0.4550 4.1690 0.6130 ;
      RECT 3.6830 0.6130 4.1690 0.6630 ;
      RECT 4.5060 0.3380 4.5560 0.4050 ;
      RECT 4.1190 0.4050 4.5560 0.4550 ;
      RECT 3.0150 0.8130 3.1050 0.8630 ;
      RECT 3.0550 0.4620 3.1050 0.8130 ;
      RECT 3.0150 0.8630 3.0650 1.0830 ;
      RECT 2.9990 0.4120 3.1050 0.4620 ;
      RECT 2.2550 1.0830 3.0650 1.1330 ;
      RECT 3.0150 1.1330 3.0650 1.3540 ;
      RECT 2.2550 0.7520 2.3050 1.0830 ;
      RECT 2.2550 0.7020 2.3450 0.7520 ;
      RECT 2.2950 0.5510 2.3450 0.7020 ;
      RECT 2.2550 0.5010 2.3450 0.5510 ;
      RECT 2.2550 0.4070 2.3050 0.5010 ;
      RECT 2.4070 0.6130 2.8530 0.6630 ;
      RECT 2.4070 0.6630 2.4570 1.0040 ;
      RECT 2.4070 0.4130 2.4570 0.6130 ;
      RECT 2.6180 0.0940 3.3150 0.1440 ;
      RECT 6.4350 0.1380 6.4850 0.1700 ;
      RECT 3.5190 0.0880 6.4850 0.1380 ;
      RECT 8.3190 0.8200 8.8670 0.8700 ;
      RECT 1.6500 0.7020 1.9410 0.7280 ;
      RECT 1.6870 0.6780 1.9410 0.7020 ;
      RECT 1.3430 0.4600 1.3930 0.5020 ;
      RECT 1.0230 0.4100 1.3930 0.4600 ;
      RECT 1.0230 1.0200 1.7000 1.0700 ;
      RECT 1.6500 0.7520 1.7000 1.0200 ;
      RECT 1.6500 0.7280 1.7370 0.7520 ;
      RECT 1.6870 0.5520 1.7370 0.6780 ;
      RECT 1.3430 0.5020 1.7370 0.5520 ;
      RECT 0.8870 0.3100 1.5450 0.3600 ;
      RECT 1.4950 0.3600 1.5450 0.3920 ;
      RECT 0.8870 0.3600 0.9370 0.3920 ;
      RECT 5.6590 0.8660 5.8080 0.9160 ;
      RECT 5.7580 0.9160 5.8080 0.9670 ;
      RECT 5.7580 0.9670 5.8930 1.0170 ;
      RECT 1.9910 0.6280 2.2450 0.6520 ;
      RECT 1.9520 0.6020 2.2450 0.6280 ;
      RECT 1.9910 0.6520 2.0410 0.7780 ;
      RECT 1.9520 0.5780 2.0410 0.6020 ;
      RECT 1.9520 0.7780 2.0410 0.8280 ;
      RECT 1.9520 0.3190 2.0020 0.5780 ;
      RECT 1.9520 0.8280 2.0020 1.0760 ;
      RECT 8.6230 0.7090 9.1610 0.7590 ;
      RECT 5.2010 1.5200 8.3250 1.5700 ;
      RECT 5.1830 0.5380 5.2330 1.0200 ;
      RECT 4.6710 0.5110 5.2330 0.5380 ;
      RECT 4.6870 1.0200 5.2330 1.0700 ;
      RECT 4.6710 0.4880 5.2320 0.5110 ;
      RECT 4.4230 0.7880 4.4730 1.1200 ;
      RECT 3.3740 0.7380 4.4750 0.7880 ;
      RECT 4.2310 0.5050 4.2810 0.7380 ;
      RECT 4.6870 1.0700 4.7370 1.1200 ;
      RECT 3.9110 1.1200 4.7370 1.1700 ;
      RECT 9.2470 0.6770 9.2970 0.7680 ;
      RECT 9.2070 0.4270 9.2970 0.4620 ;
      RECT 9.2470 0.1260 9.2970 0.4270 ;
      RECT 9.2070 0.6270 9.2970 0.6770 ;
      RECT 9.2070 0.5120 9.2570 0.6270 ;
      RECT 9.0030 0.4770 9.2570 0.5120 ;
      RECT 9.0030 0.4620 9.2970 0.4770 ;
      RECT 4.4430 1.5200 5.1330 1.5700 ;
      RECT 4.8980 0.6130 5.1330 0.6630 ;
      RECT 5.4470 0.8670 5.5890 0.9170 ;
      RECT 5.4470 0.6630 5.4970 0.8670 ;
      RECT 5.4470 0.6130 5.8930 0.6630 ;
      RECT 4.5350 0.9200 4.9650 0.9700 ;
      RECT 4.9150 0.8310 4.9650 0.9200 ;
      RECT 4.5350 0.9700 4.5850 1.0340 ;
      RECT 4.5350 0.5050 4.5850 0.9200 ;
      RECT 4.2910 1.4200 5.5970 1.4700 ;
      RECT 3.3030 1.1900 3.6890 1.2400 ;
      RECT 5.8800 1.2790 6.2730 1.3290 ;
      RECT 3.2270 1.3890 3.7650 1.4390 ;
      RECT 7.3310 1.1990 8.6290 1.2490 ;
      RECT 7.9390 0.5270 8.5370 0.5770 ;
      RECT 8.4870 0.5770 8.5370 0.7700 ;
      RECT 8.4870 0.3480 8.5370 0.5270 ;
      RECT 8.1830 0.5770 8.2330 0.8870 ;
      RECT 8.1830 0.1260 8.2330 0.5270 ;
      RECT 8.6230 0.1320 8.8570 0.1820 ;
      RECT 7.8790 1.0680 8.3280 1.1180 ;
      RECT 7.8790 0.6770 7.9290 1.0680 ;
      RECT 7.8390 0.6270 7.9290 0.6770 ;
      RECT 7.8390 0.4770 7.8890 0.6270 ;
      RECT 7.8390 0.4270 7.9290 0.4770 ;
      RECT 7.8790 0.1260 7.9290 0.4270 ;
      RECT 2.9230 1.5240 3.9170 1.5740 ;
      RECT 0.7190 0.5100 1.2570 0.5600 ;
      RECT 1.1750 1.1330 1.5610 1.1830 ;
      RECT 0.7190 0.9410 0.9530 0.9910 ;
      RECT 8.8510 1.0830 9.3890 1.1330 ;
      RECT 8.3190 0.2480 9.1610 0.2980 ;
      RECT 2.8630 0.7130 2.9890 0.7630 ;
      RECT 2.8630 0.7630 2.9130 1.0330 ;
      RECT 2.9390 0.5630 2.9890 0.7130 ;
      RECT 2.8470 0.5130 2.9890 0.5630 ;
      RECT 4.8230 0.3880 5.4970 0.4380 ;
      RECT 5.4470 0.4380 5.4970 0.5630 ;
      RECT 5.4470 0.2970 5.4970 0.3880 ;
    LAYER PO ;
      RECT 9.4850 0.0660 9.5150 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 5.8370 0.0660 5.8670 0.6910 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 3.1010 0.8400 3.1310 1.6060 ;
      RECT 5.8370 0.9390 5.8670 1.6060 ;
      RECT 5.5330 0.0660 5.5630 0.6370 ;
      RECT 3.1010 0.0660 3.1310 0.6370 ;
      RECT 9.3330 0.0660 9.3630 1.6060 ;
      RECT 3.7090 0.0660 3.7390 0.6910 ;
      RECT 5.0770 0.0660 5.1070 0.6910 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 9.6370 0.0660 9.6670 1.6060 ;
      RECT 4.7730 0.8920 4.8030 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 5.5330 0.8390 5.5630 1.6060 ;
      RECT 9.7890 0.0660 9.8190 1.6060 ;
      RECT 10.2450 0.0660 10.2750 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 9.9410 0.0660 9.9710 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 10.0930 0.0660 10.1230 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 4.7730 0.0660 4.8030 0.6910 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 3.7090 0.9390 3.7390 1.6060 ;
      RECT 7.3570 0.0670 7.3870 1.6050 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 5.0770 0.8390 5.1070 1.6060 ;
    LAYER NWELL ;
      RECT 7.7120 0.4910 9.7230 1.0830 ;
      RECT -0.1150 1.5430 10.4580 1.7730 ;
      RECT -0.1150 0.6790 7.2500 1.5430 ;
      RECT 10.1830 0.6790 10.4580 1.5430 ;
  END
END RSDFFSRASX1_LVT

MACRO RSDFFSRASX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.64 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.9670 0.8420 7.8190 0.8920 ;
        RECT 6.9670 0.8920 7.0170 1.3190 ;
        RECT 7.7690 0.5120 7.8190 0.8420 ;
        RECT 7.6970 0.4520 7.8190 0.5120 ;
        RECT 6.9670 0.4020 7.8190 0.4520 ;
        RECT 6.9670 0.1490 7.0170 0.4020 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 10.6400 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 1.6470 1.1310 1.6970 1.6420 ;
        RECT 2.1030 1.1310 2.1530 1.6420 ;
        RECT 1.7990 1.1310 1.8490 1.6420 ;
        RECT 2.7110 1.2940 2.7610 1.6420 ;
        RECT 3.9670 1.2700 4.0170 1.6420 ;
        RECT 8.6790 1.4540 8.7290 1.6420 ;
        RECT 2.5390 1.2440 2.7610 1.2940 ;
        RECT 3.7580 1.2200 5.0570 1.2700 ;
        RECT 5.7510 1.4040 8.7290 1.4540 ;
        RECT 5.7510 1.2790 5.8010 1.4040 ;
        RECT 7.4230 1.0530 7.4730 1.4040 ;
        RECT 6.5110 0.9530 6.5610 1.4040 ;
        RECT 6.8150 0.9130 6.8650 1.4040 ;
        RECT 7.1190 0.9610 7.1690 1.4040 ;
    END
  END VDD

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4670 1.4650 2.6390 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 10.6400 0.0300 ;
        RECT 2.1030 0.0300 2.1530 0.3070 ;
        RECT 1.6470 0.0300 1.6970 0.4050 ;
        RECT 0.5830 0.0300 0.6330 0.5120 ;
        RECT 0.4310 0.0300 0.4810 0.4340 ;
        RECT 1.7990 0.0300 1.8490 0.4050 ;
        RECT 8.3350 0.0300 8.3850 0.4260 ;
        RECT 7.1190 0.0300 7.1690 0.3200 ;
        RECT 6.8150 0.0300 6.8650 0.4090 ;
        RECT 7.4230 0.0300 7.4730 0.2210 ;
        RECT 9.7030 0.0300 9.7530 0.4260 ;
        RECT 9.2470 0.0300 9.2970 0.1980 ;
        RECT 6.6870 0.0300 6.7370 0.2880 ;
        RECT 2.1030 0.3070 3.9770 0.3570 ;
        RECT 5.7350 0.2880 6.7370 0.3380 ;
        RECT 3.7750 0.3570 3.8250 0.5570 ;
        RECT 2.5590 0.3570 2.6090 0.5570 ;
        RECT 2.7110 0.3570 2.7610 0.5570 ;
        RECT 3.9270 0.3570 3.9770 0.5330 ;
        RECT 2.1030 0.3570 2.1530 0.4050 ;
        RECT 3.9270 0.2380 3.9770 0.3070 ;
        RECT 3.9270 0.1880 5.0570 0.2380 ;
        RECT 4.3830 0.2380 4.4330 0.3490 ;
    END
  END VSS

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.9790 0.8570 6.1350 0.9750 ;
        RECT 5.9790 0.9750 6.0290 1.0790 ;
        RECT 5.4470 1.0790 6.0290 1.1290 ;
        RECT 5.4470 1.1290 5.4970 1.3200 ;
        RECT 4.1550 1.3200 5.4970 1.3700 ;
        RECT 4.1550 1.3700 4.2050 1.4550 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.2710 0.2710 7.9690 0.3210 ;
        RECT 7.8470 0.3210 7.9690 0.3600 ;
        RECT 7.8470 0.2500 7.9690 0.2710 ;
        RECT 7.2710 0.1490 7.3210 0.2710 ;
        RECT 7.9190 0.3600 7.9690 0.9420 ;
        RECT 7.8470 0.2470 7.9610 0.2500 ;
        RECT 7.2710 0.9420 7.9690 0.9920 ;
        RECT 7.2710 0.9920 7.3210 1.3270 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.8250 0.2480 9.9350 0.3580 ;
        RECT 9.8360 0.3580 9.8860 0.5270 ;
        RECT 9.6110 0.5270 9.8860 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.7630 0.5970 4.8130 0.7050 ;
        RECT 4.6570 0.7050 4.8130 0.7310 ;
        RECT 4.6570 0.7310 5.1170 0.7810 ;
        RECT 4.6570 0.7810 4.8130 0.8150 ;
        RECT 5.0670 0.7810 5.1170 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 8.3190 0.9470 9.9370 1.0070 ;
        RECT 9.8270 0.6900 9.9370 0.9470 ;
        RECT 9.7030 0.6270 9.7530 0.9470 ;
    END
  END VDDG

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2520 1.3330 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6780 0.7250 0.7280 ;
        RECT 0.4010 0.5510 0.5110 0.6780 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 1.1610 1.0110 1.3160 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D
  OBS
    LAYER M1 ;
      RECT 3.5470 0.0880 6.4850 0.1380 ;
      RECT 3.5470 0.1380 3.5970 0.1700 ;
      RECT 1.4520 0.6020 1.6370 0.6520 ;
      RECT 0.2050 0.8410 1.5020 0.8910 ;
      RECT 1.4520 0.6520 1.5020 0.8410 ;
      RECT 0.2050 0.5260 0.2550 0.8410 ;
      RECT 0.2790 0.8910 0.3290 1.2140 ;
      RECT 0.2050 0.4760 0.3290 0.5260 ;
      RECT 0.2790 0.3160 0.3290 0.4760 ;
      RECT 0.8870 0.3100 1.5450 0.3600 ;
      RECT 1.4950 0.3600 1.5450 0.3920 ;
      RECT 0.8870 0.3600 0.9370 0.3920 ;
      RECT 1.6870 0.6780 1.9410 0.7020 ;
      RECT 1.6500 0.7020 1.9410 0.7280 ;
      RECT 1.0230 0.4100 1.3930 0.4600 ;
      RECT 1.3430 0.4600 1.3930 0.5020 ;
      RECT 1.3430 0.5020 1.7370 0.5520 ;
      RECT 1.6870 0.5520 1.7370 0.6780 ;
      RECT 1.6500 0.7280 1.7370 0.7520 ;
      RECT 1.6500 0.7520 1.7000 1.0200 ;
      RECT 1.0230 1.0200 1.7000 1.0700 ;
      RECT 0.7190 0.5100 1.2570 0.5600 ;
      RECT 3.1670 0.8540 4.0690 0.9040 ;
      RECT 3.1670 0.6130 3.2170 0.8540 ;
      RECT 3.1670 0.5630 3.3690 0.6130 ;
      RECT 3.1670 0.9040 3.2170 1.0590 ;
      RECT 3.3190 0.4070 3.3690 0.5630 ;
      RECT 3.1670 0.4130 3.2170 0.5630 ;
      RECT 3.1670 1.0590 3.5370 1.1090 ;
      RECT 3.1670 1.1090 3.2170 1.3370 ;
      RECT 1.9910 0.6280 2.2450 0.6520 ;
      RECT 1.9520 0.6020 2.2450 0.6280 ;
      RECT 1.9910 0.6520 2.0410 0.7780 ;
      RECT 1.9520 0.5780 2.0410 0.6020 ;
      RECT 1.9520 0.7780 2.0410 0.8280 ;
      RECT 1.9520 0.3190 2.0020 0.5780 ;
      RECT 1.9520 0.8280 2.0020 1.0760 ;
      RECT 2.8470 0.5130 2.9890 0.5630 ;
      RECT 2.9390 0.5630 2.9890 0.7130 ;
      RECT 2.8630 0.7130 2.9890 0.7630 ;
      RECT 2.8630 0.7630 2.9130 1.0330 ;
      RECT 2.9990 0.4120 3.1050 0.4620 ;
      RECT 3.0550 0.4620 3.1050 0.8130 ;
      RECT 3.0150 0.8130 3.1050 0.8630 ;
      RECT 3.0150 0.8630 3.0650 1.0830 ;
      RECT 2.2550 1.0830 3.0650 1.1330 ;
      RECT 3.0150 1.1330 3.0650 1.3540 ;
      RECT 2.2550 0.7520 2.3050 1.0830 ;
      RECT 2.2550 0.7020 2.3450 0.7520 ;
      RECT 2.2950 0.5510 2.3450 0.7020 ;
      RECT 2.2550 0.5010 2.3450 0.5510 ;
      RECT 2.2550 0.4070 2.3050 0.5010 ;
      RECT 2.4070 0.6130 2.8530 0.6630 ;
      RECT 2.4070 0.6630 2.4570 1.0040 ;
      RECT 2.4070 0.4130 2.4570 0.6130 ;
      RECT 2.6180 0.0940 3.3150 0.1440 ;
      RECT 5.1470 0.1880 5.7410 0.2380 ;
      RECT 5.1470 0.2380 5.1970 0.2880 ;
      RECT 4.5060 0.2880 5.1970 0.3380 ;
      RECT 4.1190 0.4550 4.1690 0.6130 ;
      RECT 3.6830 0.6130 4.1690 0.6630 ;
      RECT 4.5060 0.3380 4.5560 0.4050 ;
      RECT 4.1190 0.4050 4.5560 0.4550 ;
      RECT 4.8230 0.3880 5.4970 0.4380 ;
      RECT 5.4470 0.4380 5.4970 0.5630 ;
      RECT 5.4470 0.2970 5.4970 0.3880 ;
      RECT 5.2950 0.9670 5.5130 1.0170 ;
      RECT 5.2950 0.4380 5.3450 0.9670 ;
      RECT 5.2950 1.0170 5.3450 1.1200 ;
      RECT 5.2950 1.1700 5.3450 1.2700 ;
      RECT 4.8230 1.1200 5.3450 1.1700 ;
      RECT 6.5870 0.6420 7.1090 0.6920 ;
      RECT 5.9430 0.4500 5.9930 0.7290 ;
      RECT 5.9430 0.7290 6.3090 0.7790 ;
      RECT 6.2590 0.7790 6.3090 1.1790 ;
      RECT 6.5870 0.4500 6.6370 0.6420 ;
      RECT 5.5990 0.4000 6.6370 0.4500 ;
      RECT 5.6000 1.1790 6.3090 1.2290 ;
      RECT 5.5990 0.4500 5.6490 0.5630 ;
      RECT 5.5990 0.2970 5.6490 0.4000 ;
      RECT 5.6000 1.2290 5.6500 1.3530 ;
      RECT 4.6710 0.4880 5.2330 0.5380 ;
      RECT 5.1830 0.5380 5.2330 1.0200 ;
      RECT 4.6870 1.0200 5.2330 1.0700 ;
      RECT 4.4230 0.7880 4.4730 1.1200 ;
      RECT 3.3740 0.7380 4.4750 0.7880 ;
      RECT 4.2310 0.5050 4.2810 0.7380 ;
      RECT 4.6870 1.0700 4.7370 1.1200 ;
      RECT 3.9110 1.1200 4.7370 1.1700 ;
      RECT 4.8980 0.6130 5.1330 0.6630 ;
      RECT 5.4470 0.6130 5.8930 0.6630 ;
      RECT 5.4470 0.6630 5.4970 0.8670 ;
      RECT 5.4470 0.8670 5.5890 0.9170 ;
      RECT 4.5350 0.9200 4.9650 0.9700 ;
      RECT 4.9150 0.8310 4.9650 0.9200 ;
      RECT 4.5350 0.9700 4.5850 1.0340 ;
      RECT 4.5350 0.5050 4.5850 0.9200 ;
      RECT 7.1790 0.6130 7.7170 0.6630 ;
      RECT 7.1790 0.6630 7.2290 0.7420 ;
      RECT 6.3590 0.7420 7.2290 0.7920 ;
      RECT 6.3590 0.7920 6.4090 1.3010 ;
      RECT 6.3590 0.5500 6.4090 0.7420 ;
      RECT 6.1310 0.5000 6.4090 0.5500 ;
      RECT 6.1310 0.5500 6.1810 0.6790 ;
      RECT 6.6630 0.7920 6.7130 1.3010 ;
      RECT 8.2430 0.5270 8.8410 0.5770 ;
      RECT 8.7910 0.5770 8.8410 0.7700 ;
      RECT 8.7910 0.3480 8.8410 0.5270 ;
      RECT 8.4870 0.5770 8.5370 0.8870 ;
      RECT 8.4870 0.1260 8.5370 0.5270 ;
      RECT 8.1820 1.0670 8.6310 1.1170 ;
      RECT 8.1830 0.6770 8.2330 1.0670 ;
      RECT 8.1430 0.6270 8.2330 0.6770 ;
      RECT 8.1430 0.4770 8.1930 0.6270 ;
      RECT 8.1430 0.4270 8.2330 0.4770 ;
      RECT 8.1830 0.1260 8.2330 0.4270 ;
      RECT 8.6230 0.2480 9.4650 0.2980 ;
      RECT 9.5510 0.6770 9.6010 0.7680 ;
      RECT 9.5110 0.4270 9.6010 0.4620 ;
      RECT 9.5510 0.1260 9.6010 0.4270 ;
      RECT 9.5110 0.6270 9.6010 0.6770 ;
      RECT 9.5110 0.5120 9.5610 0.6270 ;
      RECT 9.3070 0.4770 9.5610 0.5120 ;
      RECT 9.3070 0.4620 9.6010 0.4770 ;
      RECT 8.9270 0.1320 9.1610 0.1820 ;
      RECT 0.7190 0.9410 0.9530 0.9910 ;
      RECT 1.1750 1.1330 1.5610 1.1830 ;
      RECT 3.3030 1.1900 3.6890 1.2400 ;
      RECT 3.2270 1.3890 3.7650 1.4390 ;
      RECT 3.6830 0.9680 4.2630 1.0180 ;
      RECT 4.2130 0.9080 4.2630 0.9680 ;
      RECT 4.2130 0.8580 4.3730 0.9080 ;
      RECT 2.9230 1.5240 3.9170 1.5740 ;
      RECT 5.7580 0.9670 5.8930 1.0170 ;
      RECT 5.7580 0.9160 5.8080 0.9670 ;
      RECT 5.6590 0.8660 5.8080 0.9160 ;
      RECT 4.4430 1.5200 5.1330 1.5700 ;
      RECT 4.2910 1.4200 5.5970 1.4700 ;
      RECT 5.8800 1.2790 6.2730 1.3290 ;
      RECT 7.6350 1.1990 8.9330 1.2490 ;
      RECT 8.6230 0.8200 9.1710 0.8700 ;
      RECT 8.9270 0.7090 9.4650 0.7590 ;
      RECT 9.1550 1.0670 9.6970 1.1170 ;
      RECT 5.2010 1.5200 8.6290 1.5700 ;
      RECT 6.4350 0.1380 6.4850 0.1700 ;
    LAYER PO ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 3.7090 0.9390 3.7390 1.6060 ;
      RECT 7.6610 0.0670 7.6910 1.6050 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 9.3330 0.0660 9.3630 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 5.0770 0.8390 5.1070 1.6060 ;
      RECT 9.7890 0.0660 9.8190 1.6060 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 9.4850 0.0660 9.5150 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 5.8370 0.0660 5.8670 0.6910 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 3.1010 0.8400 3.1310 1.6060 ;
      RECT 5.8370 0.9390 5.8670 1.6060 ;
      RECT 5.5330 0.0660 5.5630 0.6370 ;
      RECT 3.1010 0.0660 3.1310 0.6370 ;
      RECT 3.7090 0.0660 3.7390 0.6910 ;
      RECT 9.6370 0.0660 9.6670 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 5.0770 0.0660 5.1070 0.6910 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 9.9410 0.0660 9.9710 1.6060 ;
      RECT 4.7730 0.8920 4.8030 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 5.5330 0.8390 5.5630 1.6060 ;
      RECT 10.0930 0.0660 10.1230 1.6060 ;
      RECT 10.5490 0.0660 10.5790 1.6060 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 10.2450 0.0660 10.2750 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 10.3970 0.0660 10.4270 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 4.7730 0.0660 4.8030 0.6910 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
    LAYER NWELL ;
      RECT 8.0160 0.4910 10.0270 1.0830 ;
      RECT -0.1150 1.5430 10.7620 1.7730 ;
      RECT -0.1150 0.6790 7.5540 1.5430 ;
      RECT 10.4870 0.6790 10.7620 1.5430 ;
  END
END RSDFFSRASX2_LVT

MACRO RSDFFSRSSRX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.88 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 0.1070 0.5110 0.2010 ;
        RECT 0.4010 0.2010 0.7250 0.2510 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END RSTB

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7010 0.4210 0.7510 ;
        RECT 0.2490 0.7510 0.3590 0.8250 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SETB

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9470 0.5630 1.1190 0.6730 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0290 0.8280 2.1830 0.9670 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2510 1.4160 1.6370 1.4660 ;
        RECT 1.3130 1.3230 1.4230 1.4160 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.0650 0.2480 9.1750 0.3580 ;
        RECT 9.0760 0.3580 9.1260 0.5030 ;
        RECT 8.8510 0.5030 9.1260 0.5530 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.3520 0.7680 4.8130 0.8180 ;
        RECT 4.3520 0.7050 4.5090 0.7680 ;
        RECT 4.7630 0.8180 4.8130 0.9700 ;
        RECT 4.4590 0.6340 4.5090 0.7050 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3150 1.4650 2.4870 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 9.8800 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.3550 ;
        RECT 2.3310 0.0300 2.3810 0.2740 ;
        RECT 6.5110 0.0300 6.5610 0.2410 ;
        RECT 8.9430 0.0300 8.9930 0.4260 ;
        RECT 8.4870 0.0300 8.5370 0.1980 ;
        RECT 1.1910 0.0300 1.2410 0.3590 ;
        RECT 2.1030 0.0300 2.1530 0.3740 ;
        RECT 7.5750 0.0300 7.6250 0.4260 ;
        RECT 6.2310 0.0300 6.2810 0.3340 ;
        RECT 0.2790 0.3550 0.6330 0.4050 ;
        RECT 2.3310 0.2740 3.8250 0.3240 ;
        RECT 5.4310 0.3340 6.2810 0.3840 ;
        RECT 0.5830 0.4050 0.6330 0.5290 ;
        RECT 0.2790 0.4050 0.3290 0.5130 ;
        RECT 3.6230 0.3240 3.6730 0.5570 ;
        RECT 3.7750 0.3240 3.8250 0.3470 ;
        RECT 2.5590 0.3240 2.6090 0.5570 ;
        RECT 2.4070 0.3240 2.4570 0.5570 ;
        RECT 3.7750 0.2650 3.8250 0.2740 ;
        RECT 3.7750 0.2150 4.7530 0.2650 ;
        RECT 4.0790 0.2650 4.1290 0.3920 ;
    END
  END VSS

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.3590 0.1570 6.4090 0.4010 ;
        RECT 6.3590 0.4010 7.0590 0.4510 ;
        RECT 6.9370 0.4510 7.0590 0.5380 ;
        RECT 7.0090 0.5380 7.0590 0.8590 ;
        RECT 6.3590 0.8590 7.0590 0.9090 ;
        RECT 6.3590 0.9090 6.4090 1.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 9.8800 1.7020 ;
        RECT 2.1030 1.3020 2.1530 1.6420 ;
        RECT 3.8150 1.2700 3.8650 1.6420 ;
        RECT 0.2790 1.3460 0.3290 1.6420 ;
        RECT 1.1510 1.2850 1.2010 1.6420 ;
        RECT 7.9190 1.4540 7.9690 1.6420 ;
        RECT 2.5590 1.3880 2.6090 1.6420 ;
        RECT 3.6060 1.2200 4.7530 1.2700 ;
        RECT 0.2790 1.2960 0.6330 1.3460 ;
        RECT 1.1510 1.2350 1.2570 1.2850 ;
        RECT 5.4470 1.4040 7.9690 1.4540 ;
        RECT 2.3870 1.3380 2.6090 1.3880 ;
        RECT 0.2790 0.9300 0.3290 1.2960 ;
        RECT 0.5830 0.9800 0.6330 1.2960 ;
        RECT 5.4470 1.2790 5.4970 1.4040 ;
        RECT 6.5110 0.9590 6.5610 1.4040 ;
        RECT 6.0550 0.9530 6.1050 1.4040 ;
    END
  END VDD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.6630 0.9690 7.1970 1.0190 ;
        RECT 7.1470 0.3510 7.1970 0.9690 ;
        RECT 6.6630 1.0190 6.8950 1.1290 ;
        RECT 6.6470 0.3010 7.1970 0.3510 ;
        RECT 6.6630 1.1290 6.7130 1.3270 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 7.5590 0.9420 9.1770 1.0020 ;
        RECT 9.0670 0.6900 9.1770 0.9420 ;
        RECT 8.9430 0.6270 8.9930 0.9420 ;
    END
  END VDDG
  OBS
    LAYER M1 ;
      RECT 3.9690 0.8580 4.0690 0.9080 ;
      RECT 2.7110 0.7130 2.8370 0.7630 ;
      RECT 2.7110 0.7630 2.7610 1.0330 ;
      RECT 2.7870 0.5630 2.8370 0.7130 ;
      RECT 2.6950 0.5130 2.8370 0.5630 ;
      RECT 3.0150 0.8670 3.9170 0.9170 ;
      RECT 3.0150 0.9170 3.0650 1.0590 ;
      RECT 3.0150 0.6130 3.0650 0.8670 ;
      RECT 3.0150 1.0590 3.3850 1.1090 ;
      RECT 3.0150 0.5630 3.2170 0.6130 ;
      RECT 3.0150 1.1090 3.0650 1.3370 ;
      RECT 3.1670 0.4070 3.2170 0.5630 ;
      RECT 3.0150 0.4130 3.0650 0.5630 ;
      RECT 4.5190 0.4210 5.1930 0.4710 ;
      RECT 5.1430 0.4710 5.1930 0.5950 ;
      RECT 5.1430 0.3290 5.1930 0.4210 ;
      RECT 4.9910 0.4710 5.0410 0.9670 ;
      RECT 4.9910 0.9670 5.2090 1.0170 ;
      RECT 4.9910 1.0170 5.0410 1.1200 ;
      RECT 4.9910 1.1700 5.0410 1.2700 ;
      RECT 4.5190 1.1200 5.0410 1.1700 ;
      RECT 4.8790 0.5710 4.9290 1.0200 ;
      RECT 4.3670 0.5220 4.9290 0.5710 ;
      RECT 4.3670 0.5210 4.9280 0.5220 ;
      RECT 4.3830 1.0200 4.9290 1.0700 ;
      RECT 4.1190 0.8080 4.1690 1.1200 ;
      RECT 3.2220 0.7580 4.1690 0.8080 ;
      RECT 3.9270 0.5420 3.9770 0.7580 ;
      RECT 4.3830 1.0700 4.4330 1.1200 ;
      RECT 3.9060 1.1200 4.4330 1.1700 ;
      RECT 2.2550 0.6130 2.7010 0.6630 ;
      RECT 2.2550 0.6630 2.3050 1.0040 ;
      RECT 2.2550 0.4130 2.3050 0.6130 ;
      RECT 4.8430 0.2280 5.4370 0.2780 ;
      RECT 3.7950 0.4920 3.8450 0.6580 ;
      RECT 3.5310 0.6580 3.8450 0.7080 ;
      RECT 4.8430 0.2780 4.8930 0.3210 ;
      RECT 4.2020 0.3210 4.8930 0.3710 ;
      RECT 4.2020 0.3710 4.2520 0.4420 ;
      RECT 3.7950 0.4420 4.2520 0.4920 ;
      RECT 2.4660 0.0940 3.1630 0.1440 ;
      RECT 5.4870 0.1650 5.5370 0.2000 ;
      RECT 5.4870 0.2000 6.0290 0.2500 ;
      RECT 5.9790 0.1040 6.0290 0.2000 ;
      RECT 3.3790 0.1150 5.5370 0.1650 ;
      RECT 8.7510 0.3890 8.8410 0.4390 ;
      RECT 8.7910 0.1260 8.8410 0.3890 ;
      RECT 8.7510 0.6270 8.8410 0.6770 ;
      RECT 8.7910 0.6770 8.8410 0.7680 ;
      RECT 8.7510 0.4390 8.8010 0.4620 ;
      RECT 8.5470 0.4620 8.8010 0.5120 ;
      RECT 8.7510 0.5120 8.8010 0.6270 ;
      RECT 7.4230 1.0820 7.8720 1.1320 ;
      RECT 7.4230 0.6770 7.4730 1.0820 ;
      RECT 7.3830 0.6270 7.4730 0.6770 ;
      RECT 7.3830 0.4770 7.4330 0.6270 ;
      RECT 7.3830 0.4270 7.4730 0.4770 ;
      RECT 7.4230 0.1260 7.4730 0.4270 ;
      RECT 7.4830 0.5270 8.0810 0.5770 ;
      RECT 7.7270 0.5770 7.7770 0.8690 ;
      RECT 7.7270 0.1260 7.7770 0.5270 ;
      RECT 8.0310 0.5770 8.0810 0.7700 ;
      RECT 8.0310 0.3480 8.0810 0.5270 ;
      RECT 6.5350 0.6130 6.9570 0.6630 ;
      RECT 6.5350 0.6630 6.5850 0.7590 ;
      RECT 5.8110 0.7590 6.5850 0.7620 ;
      RECT 5.9030 0.7620 6.5850 0.8090 ;
      RECT 5.8110 0.7120 5.9530 0.7590 ;
      RECT 5.9030 0.8090 5.9530 1.3010 ;
      RECT 5.9030 0.5340 5.9530 0.7120 ;
      RECT 6.2070 0.8090 6.2570 1.3010 ;
      RECT 7.8630 0.2480 8.7050 0.2980 ;
      RECT 3.1510 1.1900 3.5370 1.2400 ;
      RECT 6.8750 1.1990 8.1730 1.2490 ;
      RECT 3.9870 1.4200 5.2930 1.4700 ;
      RECT 4.2310 0.9200 4.6610 0.9700 ;
      RECT 4.6110 0.8880 4.6610 0.9200 ;
      RECT 4.2310 0.9700 4.2810 1.0340 ;
      RECT 4.2310 0.5420 4.2810 0.9200 ;
      RECT 2.8470 0.4120 2.9530 0.4620 ;
      RECT 2.9030 0.4620 2.9530 0.8130 ;
      RECT 2.8630 0.8130 2.9530 0.8630 ;
      RECT 2.8630 0.8630 2.9130 1.2020 ;
      RECT 2.8630 1.2520 2.9130 1.3540 ;
      RECT 1.6470 1.2020 2.9130 1.2520 ;
      RECT 1.6470 0.3490 1.6970 1.2020 ;
      RECT 5.4540 0.9670 5.5890 1.0170 ;
      RECT 5.4540 0.9160 5.5040 0.9670 ;
      RECT 5.3550 0.8660 5.5040 0.9160 ;
      RECT 2.7710 1.5240 3.7650 1.5740 ;
      RECT 8.1670 0.7090 8.7050 0.7590 ;
      RECT 7.8630 0.8200 8.4110 0.8700 ;
      RECT 8.1670 0.1320 8.4010 0.1820 ;
      RECT 8.3950 1.0840 8.9330 1.1340 ;
      RECT 5.6590 0.0940 5.8930 0.1440 ;
      RECT 5.1430 0.7060 5.5890 0.7560 ;
      RECT 5.1430 0.7560 5.1930 0.8670 ;
      RECT 5.1430 0.8670 5.2850 0.9170 ;
      RECT 4.5940 0.6680 4.8290 0.7180 ;
      RECT 1.2910 0.3190 1.3930 0.3690 ;
      RECT 1.3430 0.3690 1.3930 1.0020 ;
      RECT 1.2910 0.1510 1.3410 0.3190 ;
      RECT 1.2910 0.1010 1.9410 0.1510 ;
      RECT 0.8710 0.4430 1.2500 0.4930 ;
      RECT 1.2000 0.4930 1.2500 1.0520 ;
      RECT 0.8870 1.0520 1.5450 1.1020 ;
      RECT 1.4950 1.1020 1.5450 1.2520 ;
      RECT 1.4950 0.3490 1.5450 1.0520 ;
      RECT 0.8870 1.1020 0.9370 1.2460 ;
      RECT 0.8870 0.9800 0.9370 1.0520 ;
      RECT 0.7000 0.5730 0.8770 0.6230 ;
      RECT 0.7000 0.6230 0.7500 0.8440 ;
      RECT 0.4310 0.8440 0.7500 0.8940 ;
      RECT 0.4310 0.8940 0.4810 1.2460 ;
      RECT 0.4310 0.4550 0.4810 0.6010 ;
      RECT 0.4710 0.6510 0.5210 0.8440 ;
      RECT 0.4310 0.6010 0.5210 0.6510 ;
      RECT 1.4030 0.2040 1.7890 0.2540 ;
      RECT 0.7190 0.3010 1.1050 0.3510 ;
      RECT 1.7990 0.3490 2.0010 0.3990 ;
      RECT 1.9510 0.3990 2.0010 0.5370 ;
      RECT 1.7990 1.0240 2.0170 1.0740 ;
      RECT 1.7990 0.3990 1.8490 1.0240 ;
      RECT 0.4910 1.4160 0.8770 1.4660 ;
      RECT 0.7350 1.3160 1.0890 1.3660 ;
      RECT 0.7350 0.9800 0.7850 1.3160 ;
      RECT 1.0390 1.1920 1.0890 1.3160 ;
      RECT 1.7070 1.4160 1.9460 1.4660 ;
      RECT 3.0750 1.3890 3.6130 1.4390 ;
      RECT 4.1390 1.5200 4.8290 1.5700 ;
      RECT 4.8970 1.5200 7.8690 1.5700 ;
      RECT 6.1310 0.6580 6.4850 0.7080 ;
      RECT 6.4350 0.6230 6.4850 0.6580 ;
      RECT 5.2950 0.4840 5.3450 0.5950 ;
      RECT 5.2950 0.3290 5.3450 0.4340 ;
      RECT 5.2960 1.2290 5.3460 1.3530 ;
      RECT 5.6660 0.4840 5.7160 0.8140 ;
      RECT 5.6660 0.8140 5.8530 0.8640 ;
      RECT 5.8030 0.8640 5.8530 1.1790 ;
      RECT 5.2960 1.1790 5.8530 1.2290 ;
      RECT 6.1310 0.4840 6.1810 0.6580 ;
      RECT 5.2950 0.4340 6.1810 0.4840 ;
      RECT 3.5310 0.9680 4.0190 1.0180 ;
      RECT 3.9690 0.9080 4.0190 0.9680 ;
    LAYER PO ;
      RECT 0.8210 0.8700 0.8510 1.6060 ;
      RECT 1.7330 0.8700 1.7630 1.6060 ;
      RECT 0.8210 0.0760 0.8510 0.6510 ;
      RECT 1.7330 0.0760 1.7630 0.6000 ;
      RECT 1.5810 0.0760 1.6110 0.6000 ;
      RECT 0.6690 0.0760 0.6990 0.5970 ;
      RECT 4.7730 0.0660 4.8030 0.7220 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 2.9490 0.8400 2.9790 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 2.9490 0.0660 2.9790 0.6370 ;
      RECT 3.5570 0.9390 3.5870 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 4.4690 0.0660 4.4990 0.7080 ;
      RECT 5.5330 0.9390 5.5630 1.6060 ;
      RECT 4.4690 0.8920 4.4990 1.6060 ;
      RECT 4.7730 0.9010 4.8030 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 3.7090 0.0660 3.7390 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 5.2290 0.0660 5.2590 0.6740 ;
      RECT 5.5330 0.0660 5.5630 0.7770 ;
      RECT 5.2290 0.8390 5.2590 1.6060 ;
      RECT 6.9010 0.0670 6.9310 1.6050 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 3.5570 0.0660 3.5870 0.7180 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 9.6370 0.0660 9.6670 1.6060 ;
      RECT 9.4850 0.0660 9.5150 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 9.7890 0.0660 9.8190 1.6060 ;
      RECT 9.3330 0.0660 9.3630 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 1.4290 0.0760 1.4590 1.6060 ;
      RECT 0.9730 0.0760 1.0030 1.6060 ;
      RECT 2.0370 0.0760 2.0670 1.6060 ;
      RECT 1.8850 0.0760 1.9150 1.6060 ;
      RECT 1.2770 0.0760 1.3070 1.6060 ;
      RECT 2.1890 0.0760 2.2190 1.6060 ;
      RECT 0.5170 0.0760 0.5470 1.6060 ;
      RECT 1.1250 0.0760 1.1550 1.6060 ;
      RECT 0.3650 0.0760 0.3950 1.6060 ;
      RECT 0.6690 0.8160 0.6990 1.6060 ;
      RECT 1.5810 0.8700 1.6110 1.6060 ;
    LAYER NWELL ;
      RECT -0.1150 1.5430 10.0020 1.7730 ;
      RECT -0.1150 0.6790 6.7940 1.5430 ;
      RECT 9.7270 0.6790 10.0020 1.5430 ;
      RECT 7.2560 0.4910 9.2670 1.0830 ;
  END
END RSDFFSRSSRX1_LVT

MACRO RSDFFSRSSRX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.184 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 0.1070 0.5110 0.2010 ;
        RECT 0.4010 0.2010 0.7250 0.2510 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END RSTB

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7010 0.4210 0.7510 ;
        RECT 0.2490 0.7510 0.3590 0.8250 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SETB

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9470 0.5630 1.1190 0.6730 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0290 0.8280 2.1830 0.9670 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2510 1.4160 1.6370 1.4660 ;
        RECT 1.3130 1.3230 1.4230 1.4160 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.8150 0.1490 6.8650 0.2710 ;
        RECT 6.8150 0.2710 7.5130 0.3210 ;
        RECT 7.3920 0.3210 7.5130 0.3600 ;
        RECT 7.3920 0.2500 7.5130 0.2710 ;
        RECT 7.4630 0.3600 7.5130 0.9420 ;
        RECT 7.3920 0.2450 7.5050 0.2500 ;
        RECT 6.8150 0.9420 7.5130 0.9920 ;
        RECT 6.8150 0.9920 6.8650 1.3270 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.5110 0.1490 6.5610 0.4020 ;
        RECT 6.5110 0.4020 7.3630 0.4520 ;
        RECT 7.2410 0.4520 7.3630 0.5120 ;
        RECT 7.3130 0.5120 7.3630 0.8420 ;
        RECT 6.5110 0.8420 7.3630 0.8920 ;
        RECT 6.5110 0.8920 6.5610 1.3190 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.3690 0.2490 9.4790 0.3590 ;
        RECT 9.3800 0.3590 9.4300 0.5270 ;
        RECT 9.1550 0.5270 9.4300 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.3530 0.7310 4.8130 0.7810 ;
        RECT 4.3530 0.7050 4.5090 0.7310 ;
        RECT 4.3530 0.7810 4.5090 0.8150 ;
        RECT 4.7630 0.7810 4.8130 0.9330 ;
        RECT 4.4590 0.5970 4.5090 0.7050 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3150 1.4650 2.4870 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 10.1840 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.3550 ;
        RECT 2.3310 0.0300 2.3810 0.2740 ;
        RECT 9.2470 0.0300 9.2970 0.4260 ;
        RECT 6.6630 0.0300 6.7130 0.3200 ;
        RECT 6.9670 0.0300 7.0170 0.2210 ;
        RECT 8.7910 0.0300 8.8410 0.1980 ;
        RECT 1.1910 0.0300 1.2410 0.3590 ;
        RECT 2.1030 0.0300 2.1530 0.3740 ;
        RECT 6.3590 0.0300 6.4090 0.4090 ;
        RECT 7.8790 0.0300 7.9290 0.4260 ;
        RECT 6.2310 0.0300 6.2810 0.3000 ;
        RECT 0.2790 0.3550 0.6330 0.4050 ;
        RECT 2.3310 0.2740 3.8250 0.3240 ;
        RECT 5.4310 0.3000 6.2810 0.3500 ;
        RECT 0.5830 0.4050 0.6330 0.5290 ;
        RECT 0.2790 0.4050 0.3290 0.5130 ;
        RECT 3.6230 0.3240 3.6730 0.5570 ;
        RECT 3.7750 0.3240 3.8250 0.3470 ;
        RECT 2.5590 0.3240 2.6090 0.5570 ;
        RECT 2.4070 0.3240 2.4570 0.5570 ;
        RECT 3.7750 0.2380 3.8250 0.2740 ;
        RECT 3.7750 0.1880 4.7530 0.2380 ;
        RECT 4.0790 0.2380 4.1290 0.3490 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 10.1840 1.7020 ;
        RECT 2.1030 1.3020 2.1530 1.6420 ;
        RECT 3.8150 1.2700 3.8650 1.6420 ;
        RECT 0.2790 1.3460 0.3290 1.6420 ;
        RECT 1.1510 1.2850 1.2010 1.6420 ;
        RECT 8.2230 1.4540 8.2730 1.6420 ;
        RECT 2.5590 1.3880 2.6090 1.6420 ;
        RECT 3.6060 1.2200 4.7530 1.2700 ;
        RECT 0.2790 1.2960 0.6330 1.3460 ;
        RECT 1.1510 1.2350 1.2570 1.2850 ;
        RECT 5.4470 1.4040 8.2730 1.4540 ;
        RECT 2.3870 1.3380 2.6090 1.3880 ;
        RECT 0.2790 0.9300 0.3290 1.2960 ;
        RECT 0.5830 0.9800 0.6330 1.2960 ;
        RECT 5.4470 1.2790 5.4970 1.4040 ;
        RECT 6.6630 0.9610 6.7130 1.4040 ;
        RECT 6.9670 1.0530 7.0170 1.4040 ;
        RECT 6.3590 0.9130 6.4090 1.4040 ;
        RECT 6.0550 0.9530 6.1050 1.4040 ;
    END
  END VDD

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 7.8630 0.9470 9.4810 1.0070 ;
        RECT 9.3710 0.6900 9.4810 0.9470 ;
        RECT 9.2470 0.6270 9.2970 0.9470 ;
    END
  END VDDG
  OBS
    LAYER M1 ;
      RECT 5.8030 0.7790 5.8530 1.1790 ;
      RECT 5.2960 1.1790 5.8530 1.2290 ;
      RECT 6.1310 0.4500 6.1810 0.6420 ;
      RECT 5.2950 0.4000 6.1810 0.4500 ;
      RECT 3.5310 0.9680 4.0190 1.0180 ;
      RECT 3.9690 0.9080 4.0190 0.9680 ;
      RECT 3.9690 0.8580 4.0690 0.9080 ;
      RECT 2.7110 0.7130 2.8370 0.7630 ;
      RECT 2.7110 0.7630 2.7610 1.0330 ;
      RECT 2.7870 0.5630 2.8370 0.7130 ;
      RECT 2.6950 0.5130 2.8370 0.5630 ;
      RECT 3.0150 0.8540 3.9170 0.9040 ;
      RECT 3.0150 0.9040 3.0650 1.0590 ;
      RECT 3.0150 0.6130 3.0650 0.8540 ;
      RECT 3.0150 1.0590 3.3850 1.1090 ;
      RECT 3.0150 0.5630 3.2170 0.6130 ;
      RECT 3.0150 1.1090 3.0650 1.3370 ;
      RECT 3.1670 0.4070 3.2170 0.5630 ;
      RECT 3.0150 0.4130 3.0650 0.5630 ;
      RECT 4.9910 1.0170 5.0410 1.1200 ;
      RECT 4.9910 0.9670 5.2090 1.0170 ;
      RECT 4.9910 1.1700 5.0410 1.2700 ;
      RECT 4.9910 0.4380 5.0410 0.9670 ;
      RECT 4.5190 0.3880 5.1930 0.4380 ;
      RECT 5.1430 0.4380 5.1930 0.5630 ;
      RECT 5.1430 0.2970 5.1930 0.3880 ;
      RECT 4.5190 1.1200 5.0410 1.1700 ;
      RECT 2.2550 0.6130 2.7010 0.6630 ;
      RECT 2.2550 0.6630 2.3050 1.0040 ;
      RECT 2.2550 0.4130 2.3050 0.6130 ;
      RECT 4.8430 0.1880 5.4370 0.2380 ;
      RECT 3.7950 0.4550 3.8450 0.6130 ;
      RECT 3.5310 0.6130 3.8450 0.6630 ;
      RECT 4.8430 0.2380 4.8930 0.2880 ;
      RECT 4.2020 0.3380 4.2520 0.4050 ;
      RECT 3.7950 0.4050 4.2520 0.4550 ;
      RECT 4.2020 0.2880 4.8930 0.3380 ;
      RECT 2.4660 0.0940 3.1630 0.1440 ;
      RECT 5.4870 0.1380 5.5370 0.2000 ;
      RECT 5.4870 0.2000 6.0290 0.2500 ;
      RECT 5.9790 0.0880 6.0290 0.2000 ;
      RECT 3.3790 0.0880 5.5370 0.1380 ;
      RECT 9.0950 0.6770 9.1450 0.7680 ;
      RECT 9.0550 0.4270 9.1450 0.4620 ;
      RECT 9.0950 0.1260 9.1450 0.4270 ;
      RECT 9.0550 0.6270 9.1450 0.6770 ;
      RECT 9.0550 0.5120 9.1050 0.6270 ;
      RECT 8.8510 0.4770 9.1050 0.5120 ;
      RECT 8.8510 0.4620 9.1450 0.4770 ;
      RECT 7.7270 1.0710 8.1760 1.1210 ;
      RECT 7.7270 0.6770 7.7770 1.0710 ;
      RECT 7.6870 0.6270 7.7770 0.6770 ;
      RECT 7.6870 0.4770 7.7370 0.6270 ;
      RECT 7.6870 0.4270 7.7770 0.4770 ;
      RECT 7.7270 0.1260 7.7770 0.4270 ;
      RECT 7.7870 0.5270 8.3850 0.5770 ;
      RECT 8.0310 0.5770 8.0810 0.8870 ;
      RECT 8.0310 0.1260 8.0810 0.5270 ;
      RECT 8.3350 0.5770 8.3850 0.7700 ;
      RECT 8.3350 0.3480 8.3850 0.5270 ;
      RECT 6.7030 0.6130 7.2610 0.6630 ;
      RECT 5.9030 0.7920 5.9530 1.3010 ;
      RECT 5.9030 0.6780 5.9530 0.7420 ;
      RECT 5.8110 0.6280 5.9530 0.6780 ;
      RECT 5.9030 0.5000 5.9530 0.6280 ;
      RECT 6.2070 0.7920 6.2570 1.3010 ;
      RECT 6.7030 0.6630 6.7530 0.7420 ;
      RECT 5.9030 0.7420 6.7530 0.7920 ;
      RECT 8.1670 0.2480 9.0090 0.2980 ;
      RECT 7.1790 1.1990 8.4770 1.2490 ;
      RECT 3.9870 1.4200 5.2930 1.4700 ;
      RECT 4.2310 0.9200 4.6610 0.9700 ;
      RECT 4.6110 0.8310 4.6610 0.9200 ;
      RECT 4.2310 0.9700 4.2810 1.0340 ;
      RECT 4.2310 0.5050 4.2810 0.9200 ;
      RECT 2.8470 0.4120 2.9530 0.4620 ;
      RECT 2.9030 0.4620 2.9530 0.8130 ;
      RECT 2.8630 0.8130 2.9530 0.8630 ;
      RECT 2.8630 0.8630 2.9130 1.2020 ;
      RECT 2.8630 1.2520 2.9130 1.3540 ;
      RECT 1.6470 1.2020 2.9130 1.2520 ;
      RECT 1.6470 0.3490 1.6970 1.2020 ;
      RECT 4.3670 0.4880 4.9290 0.5380 ;
      RECT 4.8790 0.5380 4.9290 1.0200 ;
      RECT 4.3830 1.0200 4.9290 1.0700 ;
      RECT 4.1190 0.7880 4.1690 1.1200 ;
      RECT 3.2220 0.7380 4.1710 0.7880 ;
      RECT 3.9270 0.5050 3.9770 0.7380 ;
      RECT 4.3830 1.0700 4.4330 1.1200 ;
      RECT 3.9060 1.1200 4.4330 1.1700 ;
      RECT 5.4540 0.9670 5.5890 1.0170 ;
      RECT 5.4540 0.9160 5.5040 0.9670 ;
      RECT 5.3550 0.8660 5.5040 0.9160 ;
      RECT 2.7710 1.5240 3.7650 1.5740 ;
      RECT 8.4710 0.7090 9.0090 0.7590 ;
      RECT 8.1670 0.8200 8.7150 0.8700 ;
      RECT 8.4710 0.1320 8.7050 0.1820 ;
      RECT 8.6990 1.0760 9.2370 1.1260 ;
      RECT 5.6590 0.0940 5.8930 0.1440 ;
      RECT 5.1430 0.6130 5.5890 0.6630 ;
      RECT 5.1430 0.6630 5.1930 0.8670 ;
      RECT 5.1430 0.8670 5.2850 0.9170 ;
      RECT 4.5940 0.6130 4.8290 0.6630 ;
      RECT 1.2910 0.3190 1.3930 0.3690 ;
      RECT 1.3430 0.3690 1.3930 1.0020 ;
      RECT 1.2910 0.1510 1.3410 0.3190 ;
      RECT 1.2910 0.1010 1.9410 0.1510 ;
      RECT 0.8710 0.4430 1.2500 0.4930 ;
      RECT 1.2000 0.4930 1.2500 1.0520 ;
      RECT 0.8870 1.0520 1.5450 1.1020 ;
      RECT 1.4950 1.1020 1.5450 1.2520 ;
      RECT 1.4950 0.3490 1.5450 1.0520 ;
      RECT 0.8870 1.1020 0.9370 1.2460 ;
      RECT 0.8870 0.9800 0.9370 1.0520 ;
      RECT 0.7000 0.5730 0.8770 0.6230 ;
      RECT 0.7000 0.6230 0.7500 0.8440 ;
      RECT 0.4310 0.8440 0.7500 0.8940 ;
      RECT 0.4310 0.8940 0.4810 1.2460 ;
      RECT 0.4310 0.4550 0.4810 0.6010 ;
      RECT 0.4710 0.6510 0.5210 0.8440 ;
      RECT 0.4310 0.6010 0.5210 0.6510 ;
      RECT 1.4030 0.2040 1.7890 0.2540 ;
      RECT 0.7190 0.3010 1.1050 0.3510 ;
      RECT 1.7990 0.3490 2.0010 0.3990 ;
      RECT 1.9510 0.3990 2.0010 0.5370 ;
      RECT 1.7990 1.0240 2.0170 1.0740 ;
      RECT 1.7990 0.3990 1.8490 1.0240 ;
      RECT 0.4910 1.4160 0.8770 1.4660 ;
      RECT 0.7350 1.3160 1.0890 1.3660 ;
      RECT 0.7350 0.9800 0.7850 1.3160 ;
      RECT 1.0390 1.1920 1.0890 1.3160 ;
      RECT 1.7070 1.4160 1.9460 1.4660 ;
      RECT 3.0750 1.3890 3.6130 1.4390 ;
      RECT 4.1390 1.5200 4.8290 1.5700 ;
      RECT 4.8970 1.5200 8.1730 1.5700 ;
      RECT 3.1510 1.1900 3.5370 1.2400 ;
      RECT 6.1310 0.6420 6.6530 0.6920 ;
      RECT 5.2950 0.4500 5.3450 0.5630 ;
      RECT 5.2950 0.2970 5.3450 0.4000 ;
      RECT 5.2960 1.2290 5.3460 1.3530 ;
      RECT 5.6660 0.4500 5.7160 0.7290 ;
      RECT 5.6660 0.7290 5.8530 0.7790 ;
    LAYER PO ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 1.4290 0.0760 1.4590 1.6060 ;
      RECT 0.9730 0.0760 1.0030 1.6060 ;
      RECT 2.0370 0.0760 2.0670 1.6060 ;
      RECT 1.8850 0.0760 1.9150 1.6060 ;
      RECT 1.2770 0.0760 1.3070 1.6060 ;
      RECT 2.1890 0.0760 2.2190 1.6060 ;
      RECT 0.5170 0.0760 0.5470 1.6060 ;
      RECT 1.1250 0.0760 1.1550 1.6060 ;
      RECT 0.3650 0.0760 0.3950 1.6060 ;
      RECT 0.6690 0.8160 0.6990 1.6060 ;
      RECT 1.5810 0.8700 1.6110 1.6060 ;
      RECT 0.8210 0.8700 0.8510 1.6060 ;
      RECT 1.7330 0.8700 1.7630 1.6060 ;
      RECT 0.8210 0.0760 0.8510 0.6510 ;
      RECT 1.7330 0.0760 1.7630 0.6000 ;
      RECT 1.5810 0.0760 1.6110 0.6000 ;
      RECT 0.6690 0.0760 0.6990 0.5970 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 4.7730 0.0660 4.8030 0.6910 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 2.9490 0.8400 2.9790 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 9.4850 0.0660 9.5150 1.6060 ;
      RECT 2.9490 0.0660 2.9790 0.6370 ;
      RECT 3.5570 0.9390 3.5870 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 4.4690 0.0660 4.4990 0.6910 ;
      RECT 5.5330 0.9390 5.5630 1.6060 ;
      RECT 4.4690 0.8920 4.4990 1.6060 ;
      RECT 4.7730 0.8390 4.8030 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 3.7090 0.0660 3.7390 1.6060 ;
      RECT 3.5570 0.0660 3.5870 0.6910 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 5.2290 0.0660 5.2590 0.6370 ;
      RECT 5.5330 0.0660 5.5630 0.6910 ;
      RECT 5.2290 0.8390 5.2590 1.6060 ;
      RECT 7.2050 0.0670 7.2350 1.6050 ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 9.3330 0.0660 9.3630 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 9.9410 0.0660 9.9710 1.6060 ;
      RECT 9.7890 0.0660 9.8190 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 10.0930 0.0660 10.1230 1.6060 ;
      RECT 9.6370 0.0660 9.6670 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
    LAYER NWELL ;
      RECT 7.5600 0.4910 9.5710 1.0830 ;
      RECT -0.1150 1.5430 10.3060 1.7730 ;
      RECT -0.1150 0.6790 7.0980 1.5430 ;
      RECT 10.0310 0.6790 10.3060 1.5430 ;
  END
END RSDFFSRSSRX2_LVT

MACRO RSDFFSRX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.728 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 9.7280 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 2.1030 1.1310 2.1530 1.6420 ;
        RECT 1.7990 1.1310 1.8490 1.6420 ;
        RECT 1.6470 1.1310 1.6970 1.6420 ;
        RECT 2.7110 1.2940 2.7610 1.6420 ;
        RECT 3.8150 1.2700 3.8650 1.6420 ;
        RECT 7.7670 1.4540 7.8170 1.6420 ;
        RECT 2.5390 1.2440 2.7610 1.2940 ;
        RECT 3.6070 1.2200 4.7530 1.2700 ;
        RECT 5.4470 1.4040 7.8170 1.4540 ;
        RECT 5.4470 1.2790 5.4970 1.4040 ;
        RECT 6.3590 0.9590 6.4090 1.4040 ;
        RECT 5.9030 0.9530 5.9530 1.4040 ;
    END
  END VDD

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.2070 0.4010 6.9070 0.4510 ;
        RECT 6.2070 0.1570 6.2570 0.4010 ;
        RECT 6.7850 0.4510 6.9070 0.5380 ;
        RECT 6.8570 0.5380 6.9070 0.8590 ;
        RECT 6.2070 0.8590 6.9070 0.9090 ;
        RECT 6.2070 0.9090 6.2570 1.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.5110 0.9690 7.0450 1.0190 ;
        RECT 6.9950 0.3510 7.0450 0.9690 ;
        RECT 6.5110 1.0190 6.7430 1.1290 ;
        RECT 6.4950 0.3010 7.0450 0.3510 ;
        RECT 6.5110 1.1290 6.5610 1.3270 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4670 1.4650 2.6390 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 9.7280 0.0300 ;
        RECT 2.1030 0.0300 2.1530 0.2570 ;
        RECT 8.7910 0.0300 8.8410 0.4260 ;
        RECT 1.6470 0.0300 1.6970 0.4050 ;
        RECT 6.3590 0.0300 6.4090 0.2410 ;
        RECT 1.7990 0.0300 1.8490 0.4050 ;
        RECT 7.4230 0.0300 7.4730 0.4260 ;
        RECT 0.5830 0.0300 0.6330 0.5120 ;
        RECT 0.4310 0.0300 0.4810 0.4340 ;
        RECT 8.3350 0.0300 8.3850 0.1980 ;
        RECT 6.0790 0.0300 6.1290 0.2830 ;
        RECT 2.1030 0.2570 3.8250 0.3070 ;
        RECT 5.4310 0.2830 6.1290 0.3330 ;
        RECT 2.5590 0.3070 2.6090 0.5570 ;
        RECT 2.7110 0.3070 2.7610 0.5570 ;
        RECT 2.1030 0.3070 2.1530 0.4050 ;
        RECT 3.7750 0.2340 3.8250 0.2570 ;
        RECT 3.7750 0.1840 4.7530 0.2340 ;
        RECT 4.0790 0.2340 4.1290 0.3490 ;
    END
  END VSS

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.9130 0.2490 9.0230 0.3590 ;
        RECT 8.9240 0.3590 8.9740 0.5050 ;
        RECT 8.6990 0.5050 8.9740 0.5550 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.3530 0.7050 4.5090 0.7310 ;
        RECT 4.3530 0.7310 4.8130 0.7810 ;
        RECT 4.4590 0.5970 4.5090 0.7050 ;
        RECT 4.3530 0.7810 4.5090 0.8150 ;
        RECT 4.7630 0.7810 4.8130 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 7.4070 0.9420 9.0250 1.0020 ;
        RECT 8.9150 0.6900 9.0250 0.9420 ;
        RECT 8.7910 0.6270 8.8410 0.9420 ;
    END
  END VDDG

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2520 1.3330 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6780 0.7250 0.7280 ;
        RECT 0.4010 0.5510 0.5110 0.6780 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 1.1610 1.0110 1.3160 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D
  OBS
    LAYER M1 ;
      RECT 3.1670 0.4340 3.3850 0.4840 ;
      RECT 3.1670 1.0990 3.3850 1.1490 ;
      RECT 3.1670 0.4080 3.2170 0.4340 ;
      RECT 3.1670 1.1490 3.2170 1.3370 ;
      RECT 1.6500 0.7020 1.9410 0.7280 ;
      RECT 1.6870 0.6780 1.9410 0.7020 ;
      RECT 1.3430 0.4600 1.3930 0.5020 ;
      RECT 1.0230 0.4100 1.3930 0.4600 ;
      RECT 1.0230 1.0200 1.7000 1.0700 ;
      RECT 1.6500 0.7520 1.7000 1.0200 ;
      RECT 1.6500 0.7280 1.7370 0.7520 ;
      RECT 1.6870 0.5520 1.7370 0.6780 ;
      RECT 1.3430 0.5020 1.7370 0.5520 ;
      RECT 0.8870 0.3100 1.5450 0.3600 ;
      RECT 1.4950 0.3600 1.5450 0.3920 ;
      RECT 0.8870 0.3600 0.9370 0.3920 ;
      RECT 5.3550 0.8660 5.5040 0.9160 ;
      RECT 5.4540 0.9160 5.5040 0.9670 ;
      RECT 5.4540 0.9670 5.5890 1.0170 ;
      RECT 6.3830 0.6130 6.8050 0.6630 ;
      RECT 5.8270 0.5670 5.8770 0.7590 ;
      RECT 6.0550 0.8090 6.1050 1.3010 ;
      RECT 5.8260 0.5170 5.9690 0.5670 ;
      RECT 6.3830 0.6630 6.4330 0.7590 ;
      RECT 5.8260 0.7590 6.4330 0.8090 ;
      RECT 1.9910 0.6280 2.2450 0.6520 ;
      RECT 1.9520 0.6020 2.2450 0.6280 ;
      RECT 1.9910 0.6520 2.0410 0.7780 ;
      RECT 1.9520 0.5780 2.0410 0.6020 ;
      RECT 1.9520 0.7780 2.0410 0.8280 ;
      RECT 1.9520 0.3190 2.0020 0.5780 ;
      RECT 1.9520 0.8280 2.0020 1.0760 ;
      RECT 2.2550 1.0830 3.0650 1.1330 ;
      RECT 3.0150 1.1330 3.0650 1.3540 ;
      RECT 3.0150 0.8630 3.0650 1.0830 ;
      RECT 3.0150 0.8130 3.1050 0.8630 ;
      RECT 3.0550 0.4620 3.1050 0.8130 ;
      RECT 2.9990 0.4120 3.1050 0.4620 ;
      RECT 2.2550 0.7520 2.3050 1.0830 ;
      RECT 2.2550 0.7020 2.3450 0.7520 ;
      RECT 2.2950 0.5510 2.3450 0.7020 ;
      RECT 2.2550 0.5010 2.3450 0.5510 ;
      RECT 2.2550 0.4070 2.3050 0.5010 ;
      RECT 8.0150 0.7090 8.5530 0.7590 ;
      RECT 3.2270 1.4240 3.6130 1.4740 ;
      RECT 2.4070 0.6130 2.8530 0.6630 ;
      RECT 2.4070 0.6630 2.4570 1.0040 ;
      RECT 2.4070 0.4130 2.4570 0.6130 ;
      RECT 4.8790 0.5340 4.9290 1.0200 ;
      RECT 4.3670 0.5070 4.9290 0.5340 ;
      RECT 4.3830 1.0200 4.9290 1.0700 ;
      RECT 4.3670 0.4840 4.9280 0.5070 ;
      RECT 4.1190 0.7880 4.1690 1.1200 ;
      RECT 3.3730 0.7380 4.1710 0.7880 ;
      RECT 3.9270 0.5050 3.9770 0.7380 ;
      RECT 4.3830 1.0700 4.4330 1.1200 ;
      RECT 3.7590 1.1200 4.4330 1.1700 ;
      RECT 8.5990 0.6270 8.6890 0.6770 ;
      RECT 8.6390 0.6770 8.6890 0.7680 ;
      RECT 8.5990 0.3770 8.6890 0.4270 ;
      RECT 8.6390 0.1260 8.6890 0.3770 ;
      RECT 8.5990 0.5120 8.6490 0.6270 ;
      RECT 8.3950 0.4620 8.6490 0.5120 ;
      RECT 8.5990 0.4270 8.6490 0.4620 ;
      RECT 4.1390 1.5200 4.8290 1.5700 ;
      RECT 4.5940 0.6130 4.8290 0.6630 ;
      RECT 5.1430 0.8670 5.2850 0.9170 ;
      RECT 5.1430 0.6630 5.1930 0.8670 ;
      RECT 5.1430 0.6130 5.5890 0.6630 ;
      RECT 4.8430 0.1780 5.4370 0.2280 ;
      RECT 4.8430 0.2280 4.8930 0.2840 ;
      RECT 4.2020 0.2840 4.8930 0.3340 ;
      RECT 3.5470 0.5240 3.5970 0.6130 ;
      RECT 3.7820 0.4550 3.8320 0.6130 ;
      RECT 3.5470 0.6130 3.8320 0.6630 ;
      RECT 4.2020 0.3340 4.2520 0.4050 ;
      RECT 3.7820 0.4050 4.2520 0.4550 ;
      RECT 4.2310 0.9200 4.6610 0.9700 ;
      RECT 4.6110 0.8310 4.6610 0.9200 ;
      RECT 4.2310 0.9700 4.2810 1.0340 ;
      RECT 4.2310 0.5050 4.2810 0.9200 ;
      RECT 3.9870 1.4200 5.2930 1.4700 ;
      RECT 6.7230 1.1990 8.0210 1.2490 ;
      RECT 2.6180 0.0940 3.3150 0.1440 ;
      RECT 7.7110 0.8200 8.2590 0.8700 ;
      RECT 8.0150 0.1320 8.2490 0.1820 ;
      RECT 7.2710 1.0870 7.7200 1.1370 ;
      RECT 7.2710 0.6770 7.3210 1.0870 ;
      RECT 7.2310 0.6270 7.3210 0.6770 ;
      RECT 7.2310 0.4770 7.2810 0.6270 ;
      RECT 7.2310 0.4270 7.3210 0.4770 ;
      RECT 7.2710 0.1260 7.3210 0.4270 ;
      RECT 2.9230 1.5240 3.7650 1.5740 ;
      RECT 7.3310 0.5270 7.9290 0.5770 ;
      RECT 7.5750 0.5770 7.6250 0.8690 ;
      RECT 7.5750 0.1260 7.6250 0.5270 ;
      RECT 7.8790 0.5770 7.9290 0.7700 ;
      RECT 7.8790 0.3480 7.9290 0.5270 ;
      RECT 5.6590 0.0960 5.8930 0.1460 ;
      RECT 0.7190 0.5100 1.2570 0.5600 ;
      RECT 1.1750 1.1330 1.5610 1.1830 ;
      RECT 0.7190 0.9410 0.9530 0.9910 ;
      RECT 8.2430 1.1000 8.7810 1.1500 ;
      RECT 7.7110 0.2480 8.5530 0.2980 ;
      RECT 4.8970 1.5200 7.7170 1.5700 ;
      RECT 2.8630 0.7130 2.9890 0.7630 ;
      RECT 2.8630 0.7630 2.9130 1.0330 ;
      RECT 2.9390 0.5630 2.9890 0.7130 ;
      RECT 2.8470 0.5130 2.9890 0.5630 ;
      RECT 4.5190 0.3840 5.1930 0.4340 ;
      RECT 5.1430 0.4340 5.1930 0.5630 ;
      RECT 5.1430 0.2970 5.1930 0.3840 ;
      RECT 4.9910 0.4340 5.0410 0.9670 ;
      RECT 4.9910 0.9670 5.2090 1.0170 ;
      RECT 4.9910 1.0170 5.0410 1.1200 ;
      RECT 4.9910 1.1700 5.0410 1.2700 ;
      RECT 4.5190 1.1200 5.0410 1.1700 ;
      RECT 3.5270 0.9680 4.0390 1.0180 ;
      RECT 3.9860 0.9080 4.0360 0.9680 ;
      RECT 3.9860 0.8580 4.0690 0.9080 ;
      RECT 1.4520 0.6020 1.6370 0.6520 ;
      RECT 0.2050 0.8410 1.5020 0.8910 ;
      RECT 1.4520 0.6520 1.5020 0.8410 ;
      RECT 0.2050 0.5260 0.2550 0.8410 ;
      RECT 0.2790 0.8910 0.3290 1.2140 ;
      RECT 0.2050 0.4760 0.3290 0.5260 ;
      RECT 0.2790 0.3160 0.3290 0.4760 ;
      RECT 5.9630 0.6320 6.3330 0.6820 ;
      RECT 6.2830 0.5970 6.3330 0.6320 ;
      RECT 5.6600 0.4500 5.7100 1.1790 ;
      RECT 5.2960 1.1790 5.8170 1.2290 ;
      RECT 6.0890 0.4500 6.1390 0.6320 ;
      RECT 5.2950 0.4000 6.1390 0.4500 ;
      RECT 5.2950 0.4500 5.3450 0.5630 ;
      RECT 5.2950 0.2970 5.3450 0.4000 ;
      RECT 5.2960 1.2290 5.3460 1.3530 ;
      RECT 3.1670 0.8540 3.9170 0.9040 ;
      RECT 3.1670 0.4840 3.2170 0.8540 ;
      RECT 3.1670 0.9040 3.2170 1.0990 ;
    LAYER PO ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.7090 0.0660 3.7390 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 3.1010 0.8400 3.1310 1.6060 ;
      RECT 5.5330 0.9390 5.5630 1.6060 ;
      RECT 5.2290 0.0660 5.2590 0.6370 ;
      RECT 3.1010 0.0660 3.1310 0.6370 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 4.7730 0.0660 4.8030 0.6910 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 4.4690 0.8920 4.4990 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 5.2290 0.8390 5.2590 1.6060 ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 9.6370 0.0660 9.6670 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 9.3330 0.0660 9.3630 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 9.4850 0.0660 9.5150 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 3.5570 0.0680 3.5870 0.6180 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 4.4690 0.0660 4.4990 0.6910 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 6.7490 0.0670 6.7790 1.6050 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 4.7730 0.8390 4.8030 1.6060 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 3.5570 0.7300 3.5870 1.6060 ;
      RECT 5.5330 0.0660 5.5630 0.6910 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
    LAYER NWELL ;
      RECT 7.1040 0.4910 9.1150 1.0830 ;
      RECT -0.1150 1.5430 9.8500 1.7730 ;
      RECT -0.1150 0.6790 6.6420 1.5430 ;
      RECT 9.5750 0.6790 9.8500 1.5430 ;
  END
END RSDFFSRX1_LVT

MACRO RSDFFSRX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.032 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.3590 0.1480 6.4090 0.4010 ;
        RECT 6.3590 0.4010 7.2120 0.4510 ;
        RECT 7.0880 0.4510 7.2120 0.5110 ;
        RECT 7.1620 0.5110 7.2120 0.8320 ;
        RECT 6.3590 0.8320 7.2120 0.8820 ;
        RECT 6.3590 0.8820 6.4090 1.3180 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.6630 0.1480 6.7130 0.2700 ;
        RECT 6.6630 0.2700 7.3620 0.3200 ;
        RECT 7.2410 0.3200 7.3620 0.3590 ;
        RECT 7.2410 0.2490 7.3620 0.2700 ;
        RECT 7.3120 0.3590 7.3620 0.9320 ;
        RECT 6.6630 0.9320 7.3620 0.9820 ;
        RECT 6.6630 0.9820 6.7130 1.3260 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 10.0320 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 2.1030 1.1310 2.1530 1.6420 ;
        RECT 1.7990 1.1310 1.8490 1.6420 ;
        RECT 1.6470 1.1310 1.6970 1.6420 ;
        RECT 8.0710 1.4540 8.1210 1.6420 ;
        RECT 2.7110 1.2940 2.7610 1.6420 ;
        RECT 3.8150 1.2700 3.8650 1.6420 ;
        RECT 5.4470 1.4040 8.1210 1.4540 ;
        RECT 2.5390 1.2440 2.7610 1.2940 ;
        RECT 3.6070 1.2200 4.7530 1.2700 ;
        RECT 5.4470 1.2790 5.4970 1.4040 ;
        RECT 5.9030 0.9530 5.9530 1.4040 ;
        RECT 6.2070 0.9120 6.2570 1.4040 ;
        RECT 6.5110 0.9600 6.5610 1.4040 ;
        RECT 6.8150 1.0520 6.8650 1.4040 ;
    END
  END VDD

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4670 1.4650 2.6390 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 10.0320 0.0300 ;
        RECT 2.1030 0.0300 2.1530 0.2570 ;
        RECT 6.8150 0.0300 6.8650 0.2200 ;
        RECT 6.5110 0.0300 6.5610 0.3190 ;
        RECT 6.2070 0.0300 6.2570 0.4080 ;
        RECT 9.0950 0.0300 9.1450 0.4260 ;
        RECT 1.6470 0.0300 1.6970 0.4050 ;
        RECT 1.7990 0.0300 1.8490 0.4050 ;
        RECT 7.7270 0.0300 7.7770 0.4260 ;
        RECT 0.5830 0.0300 0.6330 0.5120 ;
        RECT 0.4310 0.0300 0.4810 0.4340 ;
        RECT 8.6390 0.0300 8.6890 0.1980 ;
        RECT 6.0790 0.0300 6.1290 0.2830 ;
        RECT 2.1030 0.2570 3.8250 0.3070 ;
        RECT 5.4310 0.2830 6.1290 0.3330 ;
        RECT 2.5590 0.3070 2.6090 0.5570 ;
        RECT 2.7110 0.3070 2.7610 0.5570 ;
        RECT 2.1030 0.3070 2.1530 0.4050 ;
        RECT 3.7750 0.2340 3.8250 0.2570 ;
        RECT 3.7750 0.1840 4.7530 0.2340 ;
        RECT 4.0790 0.2340 4.1290 0.3490 ;
    END
  END VSS

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.2170 0.2490 9.3290 0.3590 ;
        RECT 9.2280 0.3590 9.2780 0.5270 ;
        RECT 9.0030 0.5270 9.2780 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.3530 0.7050 4.5090 0.7310 ;
        RECT 4.3530 0.7310 4.8130 0.7810 ;
        RECT 4.4590 0.5970 4.5090 0.7050 ;
        RECT 4.3530 0.7810 4.5090 0.8150 ;
        RECT 4.7630 0.7810 4.8130 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 7.7110 0.9420 9.3290 1.0020 ;
        RECT 9.2190 0.6900 9.3290 0.9420 ;
        RECT 9.0950 0.6270 9.1450 0.9420 ;
    END
  END VDDG

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2520 1.3330 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6780 0.7250 0.7280 ;
        RECT 0.4010 0.5510 0.5110 0.6780 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 1.1610 1.0110 1.3160 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D
  OBS
    LAYER M1 ;
      RECT 2.9990 0.4120 3.1050 0.4620 ;
      RECT 3.0550 0.4620 3.1050 0.8130 ;
      RECT 3.0150 0.8130 3.1050 0.8630 ;
      RECT 3.0150 0.8630 3.0650 1.0830 ;
      RECT 2.2550 1.0830 3.0650 1.1330 ;
      RECT 3.0150 1.1330 3.0650 1.3540 ;
      RECT 2.2550 0.7520 2.3050 1.0830 ;
      RECT 2.2550 0.7020 2.3450 0.7520 ;
      RECT 2.2950 0.5510 2.3450 0.7020 ;
      RECT 2.2550 0.5010 2.3450 0.5510 ;
      RECT 2.2550 0.4070 2.3050 0.5010 ;
      RECT 2.4070 0.6130 2.8530 0.6630 ;
      RECT 2.4070 0.6630 2.4570 1.0040 ;
      RECT 2.4070 0.4130 2.4570 0.6130 ;
      RECT 2.6180 0.0940 3.3150 0.1440 ;
      RECT 8.0150 0.8200 8.5630 0.8700 ;
      RECT 3.1670 0.8540 3.9170 0.9040 ;
      RECT 3.1670 0.4840 3.2170 0.8540 ;
      RECT 3.1670 0.9040 3.2170 1.0990 ;
      RECT 3.1670 0.4340 3.3850 0.4840 ;
      RECT 3.1670 1.0990 3.3850 1.1490 ;
      RECT 3.1670 0.4080 3.2170 0.4340 ;
      RECT 3.1670 1.1490 3.2170 1.3370 ;
      RECT 1.6500 0.7020 1.9410 0.7280 ;
      RECT 1.6870 0.6780 1.9410 0.7020 ;
      RECT 1.3430 0.4600 1.3930 0.5020 ;
      RECT 1.0230 0.4100 1.3930 0.4600 ;
      RECT 1.0230 1.0200 1.7000 1.0700 ;
      RECT 1.6500 0.7520 1.7000 1.0200 ;
      RECT 1.6500 0.7280 1.7370 0.7520 ;
      RECT 1.6870 0.5520 1.7370 0.6780 ;
      RECT 1.3430 0.5020 1.7370 0.5520 ;
      RECT 0.8870 0.3100 1.5450 0.3600 ;
      RECT 1.4950 0.3600 1.5450 0.3920 ;
      RECT 0.8870 0.3600 0.9370 0.3920 ;
      RECT 5.3550 0.8660 5.5040 0.9160 ;
      RECT 5.4540 0.9160 5.5040 0.9670 ;
      RECT 5.4540 0.9670 5.5890 1.0170 ;
      RECT 6.5650 0.6130 7.1100 0.6630 ;
      RECT 5.8270 0.5670 5.8770 0.7320 ;
      RECT 6.0550 0.7820 6.1050 1.3010 ;
      RECT 5.8260 0.5170 5.9690 0.5670 ;
      RECT 6.5650 0.6630 6.6150 0.7320 ;
      RECT 5.8260 0.7320 6.6150 0.7820 ;
      RECT 1.9910 0.6280 2.2450 0.6520 ;
      RECT 1.9520 0.6020 2.2450 0.6280 ;
      RECT 1.9910 0.6520 2.0410 0.7780 ;
      RECT 1.9520 0.5780 2.0410 0.6020 ;
      RECT 1.9520 0.7780 2.0410 0.8280 ;
      RECT 1.9520 0.3190 2.0020 0.5780 ;
      RECT 1.9520 0.8280 2.0020 1.0760 ;
      RECT 8.3190 0.7090 8.8570 0.7590 ;
      RECT 3.2270 1.4240 3.6130 1.4740 ;
      RECT 4.8790 0.5340 4.9290 1.0200 ;
      RECT 4.3670 0.5070 4.9290 0.5340 ;
      RECT 4.3830 1.0200 4.9290 1.0700 ;
      RECT 4.3670 0.4840 4.9280 0.5070 ;
      RECT 4.1190 0.7880 4.1690 1.1200 ;
      RECT 3.3730 0.7380 4.1710 0.7880 ;
      RECT 3.9270 0.5050 3.9770 0.7380 ;
      RECT 4.3830 1.0700 4.4330 1.1200 ;
      RECT 3.7590 1.1200 4.4330 1.1700 ;
      RECT 7.5750 1.0620 8.0240 1.1120 ;
      RECT 7.5750 0.6770 7.6250 1.0620 ;
      RECT 7.5350 0.6270 7.6250 0.6770 ;
      RECT 7.5350 0.4770 7.5850 0.6270 ;
      RECT 7.5350 0.4270 7.6250 0.4770 ;
      RECT 7.5750 0.1260 7.6250 0.4270 ;
      RECT 4.8430 0.1780 5.4370 0.2280 ;
      RECT 4.8430 0.2280 4.8930 0.2840 ;
      RECT 4.2020 0.2840 4.8930 0.3340 ;
      RECT 3.5470 0.5240 3.5970 0.6130 ;
      RECT 3.7820 0.4550 3.8320 0.6130 ;
      RECT 3.5470 0.6130 3.8320 0.6630 ;
      RECT 4.2020 0.3340 4.2520 0.4050 ;
      RECT 3.7820 0.4050 4.2520 0.4550 ;
      RECT 8.5470 1.0620 9.0850 1.1120 ;
      RECT 8.0150 0.2480 8.8570 0.2980 ;
      RECT 4.8970 1.5200 8.0210 1.5700 ;
      RECT 8.9430 0.6770 8.9930 0.7680 ;
      RECT 8.9030 0.4270 8.9930 0.4620 ;
      RECT 8.9430 0.1260 8.9930 0.4270 ;
      RECT 8.9030 0.6270 8.9930 0.6770 ;
      RECT 8.9030 0.5120 8.9530 0.6270 ;
      RECT 8.6990 0.4770 8.9530 0.5120 ;
      RECT 8.6990 0.4620 8.9930 0.4770 ;
      RECT 4.1390 1.5200 4.8290 1.5700 ;
      RECT 4.5940 0.6130 4.8290 0.6630 ;
      RECT 5.1430 0.8670 5.2850 0.9170 ;
      RECT 5.1430 0.6630 5.1930 0.8670 ;
      RECT 5.1430 0.6130 5.5890 0.6630 ;
      RECT 4.2310 0.9200 4.6610 0.9700 ;
      RECT 4.6110 0.8310 4.6610 0.9200 ;
      RECT 4.2310 0.9700 4.2810 1.0340 ;
      RECT 4.2310 0.5050 4.2810 0.9200 ;
      RECT 3.9870 1.4200 5.2930 1.4700 ;
      RECT 7.0270 1.1990 8.3250 1.2490 ;
      RECT 7.6350 0.5270 8.2330 0.5770 ;
      RECT 8.1830 0.5770 8.2330 0.7700 ;
      RECT 8.1830 0.3480 8.2330 0.5270 ;
      RECT 7.8790 0.5770 7.9290 0.8840 ;
      RECT 7.8790 0.1260 7.9290 0.5270 ;
      RECT 8.3190 0.1320 8.5530 0.1820 ;
      RECT 2.9230 1.5240 3.7650 1.5740 ;
      RECT 5.6590 0.0880 5.8930 0.1380 ;
      RECT 0.7190 0.5100 1.2570 0.5600 ;
      RECT 1.1750 1.1330 1.5610 1.1830 ;
      RECT 0.7190 0.9410 0.9530 0.9910 ;
      RECT 2.8630 0.7130 2.9890 0.7630 ;
      RECT 2.8630 0.7630 2.9130 1.0330 ;
      RECT 2.9390 0.5630 2.9890 0.7130 ;
      RECT 2.8470 0.5130 2.9890 0.5630 ;
      RECT 4.5190 0.3840 5.1930 0.4340 ;
      RECT 5.1430 0.4340 5.1930 0.5630 ;
      RECT 5.1430 0.2970 5.1930 0.3840 ;
      RECT 4.9910 0.4340 5.0410 0.9670 ;
      RECT 4.9910 0.9670 5.2090 1.0170 ;
      RECT 4.9910 1.0170 5.0410 1.1200 ;
      RECT 4.9910 1.1700 5.0410 1.2700 ;
      RECT 4.5190 1.1200 5.0410 1.1700 ;
      RECT 3.5270 0.9680 4.0390 1.0180 ;
      RECT 3.9860 0.9080 4.0360 0.9680 ;
      RECT 3.9860 0.8580 4.0690 0.9080 ;
      RECT 1.4520 0.6020 1.6370 0.6520 ;
      RECT 0.2050 0.8410 1.5020 0.8910 ;
      RECT 1.4520 0.6520 1.5020 0.8410 ;
      RECT 0.2050 0.5260 0.2550 0.8410 ;
      RECT 0.2790 0.8910 0.3290 1.2140 ;
      RECT 0.2050 0.4760 0.3290 0.5260 ;
      RECT 0.2790 0.3160 0.3290 0.4760 ;
      RECT 5.9630 0.6320 6.5010 0.6820 ;
      RECT 5.2950 0.4500 5.3450 0.5630 ;
      RECT 5.2950 0.2970 5.3450 0.4000 ;
      RECT 5.2960 1.2290 5.3460 1.3530 ;
      RECT 5.6600 0.4500 5.7100 1.1790 ;
      RECT 5.2960 1.1790 5.8170 1.2290 ;
      RECT 6.0890 0.4500 6.1390 0.6320 ;
      RECT 5.2950 0.4000 6.1390 0.4500 ;
    LAYER PO ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.7090 0.0660 3.7390 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 3.1010 0.8400 3.1310 1.6060 ;
      RECT 5.5330 0.9390 5.5630 1.6060 ;
      RECT 5.2290 0.0660 5.2590 0.6370 ;
      RECT 3.1010 0.0660 3.1310 0.6370 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 4.7730 0.0660 4.8030 0.6910 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 9.3330 0.0660 9.3630 1.6060 ;
      RECT 4.4690 0.8920 4.4990 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 5.2290 0.8390 5.2590 1.6060 ;
      RECT 9.4850 0.0660 9.5150 1.6060 ;
      RECT 9.9410 0.0660 9.9710 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 9.6370 0.0660 9.6670 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 9.7890 0.0660 9.8190 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 3.5570 0.0680 3.5870 0.6180 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 4.4690 0.0660 4.4990 0.6910 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 7.0530 0.0670 7.0830 1.6050 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 4.7730 0.8390 4.8030 1.6060 ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 3.5570 0.7300 3.5870 1.6060 ;
      RECT 5.5330 0.0660 5.5630 0.6910 ;
    LAYER NWELL ;
      RECT 7.4080 0.4910 9.4190 1.0830 ;
      RECT -0.1150 1.5430 10.1510 1.7730 ;
      RECT -0.1150 0.6790 6.9460 1.5430 ;
      RECT 9.8790 0.6790 10.1510 1.5430 ;
  END
END RSDFFSRX2_LVT

MACRO RSDFFX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.184 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 8.0150 0.9420 9.4820 1.0020 ;
        RECT 9.3720 0.6900 9.4820 0.9420 ;
    END
  END VDDG

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6780 0.7250 0.7280 ;
        RECT 0.4010 0.5510 0.5110 0.6780 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2520 1.3330 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 1.1610 1.0110 1.3160 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 10.1840 0.0300 ;
        RECT 2.4070 0.0300 2.4570 0.3070 ;
        RECT 9.0950 0.0300 9.1450 0.3120 ;
        RECT 8.7910 0.0300 8.8410 0.2020 ;
        RECT 8.0310 0.0300 8.0810 0.2060 ;
        RECT 1.7990 0.0300 1.8490 0.4050 ;
        RECT 2.2550 0.0300 2.3050 0.5570 ;
        RECT 6.9670 0.0300 7.0170 0.2410 ;
        RECT 1.6470 0.0300 1.6970 0.4050 ;
        RECT 0.5830 0.0300 0.6330 0.5120 ;
        RECT 0.4310 0.0300 0.4810 0.4340 ;
        RECT 6.7030 0.0300 6.7530 0.2830 ;
        RECT 2.4070 0.3070 3.9770 0.3570 ;
        RECT 4.8230 0.2830 6.7540 0.3330 ;
        RECT 3.9270 0.3570 3.9770 0.5770 ;
        RECT 3.3190 0.3570 3.3690 0.5580 ;
        RECT 3.4710 0.3570 3.5210 0.5580 ;
        RECT 6.6630 0.3330 6.7130 0.4430 ;
    END
  END VSS

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0730 1.4650 2.2460 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.1190 0.9690 7.6530 1.0190 ;
        RECT 7.1190 1.0190 7.3510 1.1290 ;
        RECT 7.6030 0.3510 7.6530 0.9690 ;
        RECT 7.1190 1.1290 7.1690 1.3270 ;
        RECT 7.1030 0.3010 7.6530 0.3510 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.8150 0.1570 6.8650 0.4010 ;
        RECT 6.8150 0.4010 7.5150 0.4510 ;
        RECT 7.3930 0.4510 7.5150 0.5380 ;
        RECT 7.4650 0.5380 7.5150 0.8590 ;
        RECT 6.8150 0.8590 7.5150 0.9090 ;
        RECT 6.8150 0.9090 6.8650 1.2320 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 10.1840 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 1.7990 1.1310 1.8490 1.6420 ;
        RECT 1.6470 1.1310 1.6970 1.6420 ;
        RECT 5.0310 1.3400 5.0810 1.6420 ;
        RECT 2.3670 1.3400 2.4170 1.6420 ;
        RECT 2.2370 1.2900 7.0180 1.3400 ;
        RECT 6.9670 0.9590 7.0170 1.2900 ;
        RECT 4.8390 0.9730 4.8890 1.2900 ;
    END
  END VDD

  PIN RETN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.3370 1.4080 8.7220 1.4580 ;
        RECT 8.6090 1.3130 8.7220 1.4080 ;
    END
    ANTENNAGATEAREA 0.084 ;
  END RETN
  OBS
    LAYER M1 ;
      RECT 4.5350 0.2770 4.7370 0.3270 ;
      RECT 4.5350 0.3270 4.5850 0.5560 ;
      RECT 4.6870 0.3270 4.7370 0.5130 ;
      RECT 4.6470 0.8170 4.6970 0.9740 ;
      RECT 4.6470 0.9740 4.7370 1.0240 ;
      RECT 4.6870 1.0240 4.7370 1.1900 ;
      RECT 4.5350 1.1900 4.7370 1.2400 ;
      RECT 4.5350 0.9740 4.5850 1.1900 ;
      RECT 8.6390 0.4620 8.9330 0.5120 ;
      RECT 8.6390 0.5120 8.6890 0.6350 ;
      RECT 8.6390 0.1820 8.6890 0.4620 ;
      RECT 8.3190 0.6350 8.6890 0.6850 ;
      RECT 8.3190 0.1320 8.6890 0.1820 ;
      RECT 8.1830 0.4940 8.5370 0.5440 ;
      RECT 8.4870 0.3480 8.5370 0.4940 ;
      RECT 8.1830 0.5440 8.2330 0.7600 ;
      RECT 5.2550 0.5630 5.3050 0.6270 ;
      RECT 5.0510 0.6270 5.3050 0.6770 ;
      RECT 5.2550 0.5130 6.1210 0.5630 ;
      RECT 5.2550 0.6770 5.3050 1.0670 ;
      RECT 5.2550 1.0670 6.1210 1.1170 ;
      RECT 3.3030 0.9670 3.9170 1.0170 ;
      RECT 3.1670 0.4070 3.2170 0.6190 ;
      RECT 3.4710 0.6690 3.5210 0.9670 ;
      RECT 3.1670 0.6190 3.5210 0.6690 ;
      RECT 9.2470 0.5620 9.5410 0.6120 ;
      RECT 9.3820 0.4120 9.4320 0.5620 ;
      RECT 9.2470 0.3620 9.4320 0.4120 ;
      RECT 9.2470 0.6120 9.2970 0.8320 ;
      RECT 8.0830 0.8320 9.2970 0.8820 ;
      RECT 9.2470 0.1260 9.2970 0.3620 ;
      RECT 8.0830 0.4200 8.1330 0.8320 ;
      RECT 8.0830 0.3700 8.2510 0.4200 ;
      RECT 4.9510 0.7670 5.1930 0.8170 ;
      RECT 5.1430 0.8170 5.1930 1.2400 ;
      RECT 4.9510 0.4530 5.0010 0.7670 ;
      RECT 4.8270 0.4030 5.1940 0.4530 ;
      RECT 5.1430 0.4530 5.1930 0.5770 ;
      RECT 4.8270 0.4530 4.8770 0.8670 ;
      RECT 4.7470 0.8670 4.8770 0.9170 ;
      RECT 1.9520 0.9670 3.0050 1.0170 ;
      RECT 1.9520 1.0170 2.0020 1.0760 ;
      RECT 1.9520 0.8280 2.0020 0.9670 ;
      RECT 1.9520 0.7780 2.0410 0.8280 ;
      RECT 1.9910 0.6280 2.0410 0.7780 ;
      RECT 1.9520 0.5780 2.0410 0.6280 ;
      RECT 1.9520 0.3190 2.0020 0.5780 ;
      RECT 2.5590 0.7130 2.6850 0.7630 ;
      RECT 2.5590 0.7630 2.6090 0.8670 ;
      RECT 2.6350 0.5630 2.6850 0.7130 ;
      RECT 2.5590 0.8670 2.8530 0.9170 ;
      RECT 2.5430 0.5130 2.6850 0.5630 ;
      RECT 7.3310 1.2000 8.4770 1.2500 ;
      RECT 2.4330 0.4130 2.8370 0.4630 ;
      RECT 2.7870 0.4630 2.8370 0.6800 ;
      RECT 2.4330 0.4630 2.4830 0.6130 ;
      RECT 2.1030 0.6130 2.5490 0.6630 ;
      RECT 2.1030 0.6630 2.1530 0.9120 ;
      RECT 2.1030 0.4130 2.1530 0.6130 ;
      RECT 5.3550 0.6130 6.2570 0.6630 ;
      RECT 6.2070 0.3830 6.2570 0.6130 ;
      RECT 5.5590 0.6630 5.6090 0.9670 ;
      RECT 5.5590 0.9670 6.2570 1.0170 ;
      RECT 6.2070 1.0170 6.2570 1.2400 ;
      RECT 1.6870 0.6780 1.9410 0.7020 ;
      RECT 1.6500 0.7020 1.9410 0.7280 ;
      RECT 1.0230 0.4100 1.3930 0.4600 ;
      RECT 1.3430 0.4600 1.3930 0.5020 ;
      RECT 1.3430 0.5020 1.7370 0.5520 ;
      RECT 1.6870 0.5520 1.7370 0.6780 ;
      RECT 1.6500 0.7280 1.7370 0.7520 ;
      RECT 1.6500 0.7520 1.7000 1.0200 ;
      RECT 1.0230 1.0200 1.7000 1.0700 ;
      RECT 0.8870 0.3100 1.5450 0.3600 ;
      RECT 1.4950 0.3600 1.5450 0.3920 ;
      RECT 0.8870 0.3600 0.9370 0.3920 ;
      RECT 3.7350 0.8670 4.0170 0.9170 ;
      RECT 3.9670 0.9170 4.0170 1.1270 ;
      RECT 3.0150 1.1270 4.0170 1.1770 ;
      RECT 3.0150 1.1770 3.0650 1.2400 ;
      RECT 3.0150 1.0660 3.1150 1.1270 ;
      RECT 3.0650 0.9170 3.1150 1.0660 ;
      RECT 3.0150 0.4130 3.0650 0.8670 ;
      RECT 3.0150 0.8670 3.3090 0.9170 ;
      RECT 3.7350 0.6070 3.7850 0.8670 ;
      RECT 3.7350 0.5570 3.8250 0.6070 ;
      RECT 3.7750 0.4130 3.8250 0.5570 ;
      RECT 1.1750 1.1330 1.5610 1.1830 ;
      RECT 4.4430 0.6130 4.6770 0.6630 ;
      RECT 2.4670 1.5240 4.6770 1.5740 ;
      RECT 2.6190 0.0940 4.3730 0.1440 ;
      RECT 0.7190 0.9410 0.9530 0.9910 ;
      RECT 4.2910 0.8670 4.5450 0.9170 ;
      RECT 0.7190 0.5100 1.2570 0.5600 ;
      RECT 3.8350 0.6670 4.2210 0.7170 ;
      RECT 6.7910 0.5010 7.0930 0.5510 ;
      RECT 7.0430 0.5510 7.0930 0.6790 ;
      RECT 6.7910 0.5510 6.8410 0.6130 ;
      RECT 6.4190 0.6130 6.8410 0.6630 ;
      RECT 1.4520 0.6020 1.6370 0.6520 ;
      RECT 0.2050 0.5260 0.2550 0.8410 ;
      RECT 0.2790 0.8910 0.3290 1.2140 ;
      RECT 0.2050 0.4760 0.3290 0.5260 ;
      RECT 0.2790 0.3160 0.3290 0.4760 ;
      RECT 0.2050 0.8410 1.5020 0.8910 ;
      RECT 1.4520 0.6520 1.5020 0.8410 ;
      RECT 7.8790 1.0620 8.3250 1.1120 ;
      RECT 7.8790 0.1260 7.9290 1.0620 ;
      RECT 4.4230 0.0920 6.5020 0.1420 ;
      RECT 4.4230 0.1420 4.4730 0.1940 ;
      RECT 4.3830 0.1940 4.4730 0.2440 ;
      RECT 4.3830 0.2440 4.4330 0.5130 ;
      RECT 4.2310 0.5130 4.4330 0.5630 ;
      RECT 4.2310 0.2770 4.2810 0.5130 ;
      RECT 4.2710 0.5630 4.3210 0.7670 ;
      RECT 4.1910 0.7670 4.3210 0.8170 ;
      RECT 4.1910 0.8170 4.2410 0.9670 ;
      RECT 4.1910 0.9670 4.2810 1.0170 ;
      RECT 4.2310 1.0170 4.2810 1.1900 ;
      RECT 4.2310 1.1900 4.4330 1.2400 ;
      RECT 4.3830 0.9740 4.4330 1.1900 ;
      RECT 5.5070 1.5280 9.5430 1.5780 ;
      RECT 5.6590 0.7130 5.8930 0.7630 ;
      RECT 5.9630 0.7590 7.4130 0.8090 ;
      RECT 6.8910 0.6420 6.9410 0.7590 ;
      RECT 6.5110 0.8090 6.5610 1.2400 ;
      RECT 6.3190 0.5630 6.3690 0.7590 ;
      RECT 6.3190 0.5130 6.5610 0.5630 ;
      RECT 6.5110 0.3830 6.5610 0.5130 ;
      RECT 9.0860 0.4120 9.1360 0.4620 ;
      RECT 9.0860 0.4620 9.2370 0.5120 ;
      RECT 9.0860 0.5120 9.1360 0.5890 ;
      RECT 8.9430 0.5890 9.1360 0.6390 ;
      RECT 8.9430 0.3620 9.1360 0.4120 ;
      RECT 8.9430 0.1260 8.9930 0.3620 ;
      RECT 8.9430 0.6390 8.9930 0.7750 ;
      RECT 4.6870 0.5130 4.7770 0.5630 ;
      RECT 4.7270 0.5630 4.7770 0.7670 ;
      RECT 4.6470 0.7670 4.7770 0.8170 ;
    LAYER PO ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 9.9410 0.0660 9.9710 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 5.3810 0.0660 5.4110 0.6910 ;
      RECT 9.7890 0.0660 9.8190 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 9.4850 0.0660 9.5150 1.6060 ;
      RECT 5.8370 0.0660 5.8670 0.7910 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 9.6370 0.0660 9.6670 1.6060 ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 4.4690 0.0660 4.4990 0.6910 ;
      RECT 4.0130 0.0660 4.0430 0.6370 ;
      RECT 2.7970 0.8390 2.8270 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 5.8370 0.9390 5.8670 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 3.7090 0.0660 3.7390 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 4.4690 0.8390 4.4990 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 9.3330 0.0660 9.3630 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 5.3810 0.9590 5.4110 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 7.3570 0.0670 7.3870 1.6050 ;
      RECT 3.5570 0.9390 3.5870 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 3.5570 0.0660 3.5870 0.6370 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 2.7970 0.0660 2.8270 0.6910 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 10.0930 0.0660 10.1230 1.6060 ;
      RECT 4.0130 0.9390 4.0430 1.6060 ;
    LAYER NWELL ;
      RECT -0.1160 1.5430 10.2770 1.7730 ;
      RECT -0.1160 0.6790 7.2510 1.5430 ;
      RECT 10.0190 0.6790 10.2770 1.5430 ;
      RECT 7.7130 0.4910 9.5590 1.0830 ;
  END
END RSDFFX1_LVT

MACRO RSDFFX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.488 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 8.3190 0.9420 9.7860 1.0020 ;
        RECT 9.6760 0.6900 9.7860 0.9420 ;
    END
  END VDDG

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6780 0.7250 0.7280 ;
        RECT 0.4010 0.5510 0.5110 0.6780 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2520 1.3330 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 1.1610 1.0110 1.3160 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.2710 0.2710 7.9690 0.3210 ;
        RECT 7.8490 0.3210 7.9690 0.3600 ;
        RECT 7.8490 0.2500 7.9690 0.2710 ;
        RECT 7.2710 0.1490 7.3210 0.2710 ;
        RECT 7.9190 0.3600 7.9690 0.9330 ;
        RECT 7.8490 0.2490 7.9610 0.2500 ;
        RECT 7.2710 0.9330 7.9690 0.9830 ;
        RECT 7.2710 0.9830 7.3210 1.2240 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.6970 0.4010 7.8090 0.4020 ;
        RECT 6.9670 0.4020 7.8190 0.4520 ;
        RECT 6.9670 0.1490 7.0170 0.4020 ;
        RECT 7.6970 0.4520 7.8190 0.5120 ;
        RECT 7.7690 0.5120 7.8190 0.8330 ;
        RECT 6.9670 0.8330 7.8190 0.8830 ;
        RECT 6.9670 0.8830 7.0170 1.2240 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 10.4880 0.0300 ;
        RECT 2.4070 0.0300 2.4570 0.3070 ;
        RECT 9.3990 0.0300 9.4490 0.3120 ;
        RECT 7.4230 0.0300 7.4730 0.2210 ;
        RECT 9.0950 0.0300 9.1450 0.2020 ;
        RECT 8.3350 0.0300 8.3850 0.2060 ;
        RECT 1.7990 0.0300 1.8490 0.4050 ;
        RECT 6.8150 0.0300 6.8650 0.4090 ;
        RECT 2.2550 0.0300 2.3050 0.5570 ;
        RECT 7.1190 0.0300 7.1690 0.3200 ;
        RECT 1.6470 0.0300 1.6970 0.4050 ;
        RECT 0.5830 0.0300 0.6330 0.5120 ;
        RECT 0.4310 0.0300 0.4810 0.4340 ;
        RECT 6.7030 0.0300 6.7530 0.2830 ;
        RECT 2.4070 0.3070 3.9770 0.3570 ;
        RECT 4.8230 0.2830 6.7540 0.3330 ;
        RECT 3.9270 0.3570 3.9770 0.5770 ;
        RECT 3.3190 0.3570 3.3690 0.5580 ;
        RECT 3.4710 0.3570 3.5210 0.5580 ;
        RECT 6.6630 0.3330 6.7130 0.4430 ;
    END
  END VSS

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0730 1.4650 2.2460 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 10.4880 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 1.7990 1.1310 1.8490 1.6420 ;
        RECT 1.6470 1.1310 1.6970 1.6420 ;
        RECT 2.3670 1.3400 2.4170 1.6420 ;
        RECT 5.0310 1.3400 5.0810 1.6420 ;
        RECT 2.2370 1.2900 7.4730 1.3400 ;
        RECT 7.4230 1.0530 7.4730 1.2900 ;
        RECT 7.1190 0.9610 7.1690 1.2900 ;
        RECT 6.8150 0.9130 6.8650 1.2900 ;
        RECT 4.8390 0.9730 4.8890 1.2900 ;
    END
  END VDD

  PIN RETN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.3370 1.4080 9.0260 1.4580 ;
        RECT 8.9130 1.3130 9.0260 1.4080 ;
    END
    ANTENNAGATEAREA 0.084 ;
  END RETN
  OBS
    LAYER M1 ;
      RECT 9.2470 0.1260 9.2970 0.3620 ;
      RECT 8.4870 0.4940 8.8410 0.5440 ;
      RECT 8.7910 0.3480 8.8410 0.4940 ;
      RECT 8.4870 0.5440 8.5370 0.7720 ;
      RECT 5.9630 0.7130 7.7170 0.7630 ;
      RECT 6.5110 0.7630 6.5610 1.2400 ;
      RECT 6.3190 0.5630 6.3690 0.7130 ;
      RECT 6.3190 0.5130 6.5610 0.5630 ;
      RECT 6.5110 0.3830 6.5610 0.5130 ;
      RECT 6.8910 0.6420 6.9410 0.7130 ;
      RECT 7.0430 0.6420 7.0930 0.7130 ;
      RECT 8.9430 0.4620 9.2370 0.5120 ;
      RECT 8.9430 0.5120 8.9930 0.6350 ;
      RECT 8.9430 0.1820 8.9930 0.4620 ;
      RECT 8.6230 0.6350 8.9930 0.6850 ;
      RECT 8.6230 0.1320 8.9930 0.1820 ;
      RECT 5.5070 1.5280 9.8470 1.5780 ;
      RECT 5.6590 0.7130 5.8930 0.7630 ;
      RECT 4.6870 0.5130 4.7770 0.5630 ;
      RECT 4.7270 0.5630 4.7770 0.7670 ;
      RECT 4.6470 0.7670 4.7770 0.8170 ;
      RECT 4.6870 0.3270 4.7370 0.5130 ;
      RECT 4.5350 0.2770 4.7370 0.3270 ;
      RECT 4.5350 0.3270 4.5850 0.5560 ;
      RECT 4.6470 0.8170 4.6970 0.9740 ;
      RECT 4.6470 0.9740 4.7370 1.0240 ;
      RECT 4.6870 1.0240 4.7370 1.1900 ;
      RECT 4.5350 1.1900 4.7370 1.2400 ;
      RECT 4.5350 0.9740 4.5850 1.1900 ;
      RECT 5.0510 0.6270 5.3050 0.6770 ;
      RECT 5.2550 0.5630 5.3050 0.6270 ;
      RECT 5.2550 0.6770 5.3050 1.0670 ;
      RECT 5.2550 0.5130 6.1210 0.5630 ;
      RECT 5.2550 1.0670 6.1210 1.1170 ;
      RECT 3.3030 0.9670 3.9170 1.0170 ;
      RECT 3.1670 0.4070 3.2170 0.6190 ;
      RECT 3.4710 0.6690 3.5210 0.9670 ;
      RECT 3.1670 0.6190 3.5210 0.6690 ;
      RECT 9.5510 0.5620 9.8450 0.6120 ;
      RECT 9.6860 0.4120 9.7360 0.5620 ;
      RECT 9.5510 0.3620 9.7360 0.4120 ;
      RECT 9.5510 0.6120 9.6010 0.8320 ;
      RECT 8.3870 0.8320 9.6010 0.8820 ;
      RECT 9.5510 0.1260 9.6010 0.3620 ;
      RECT 8.3870 0.4200 8.4370 0.8320 ;
      RECT 8.3870 0.3700 8.5550 0.4200 ;
      RECT 4.9510 0.7670 5.1930 0.8170 ;
      RECT 5.1430 0.8170 5.1930 1.2400 ;
      RECT 4.9510 0.4530 5.0010 0.7670 ;
      RECT 4.8270 0.4030 5.1940 0.4530 ;
      RECT 5.1430 0.4530 5.1930 0.5770 ;
      RECT 4.8270 0.4530 4.8770 0.8670 ;
      RECT 4.7470 0.8670 4.8770 0.9170 ;
      RECT 1.9520 0.9670 3.0050 1.0170 ;
      RECT 1.9520 1.0170 2.0020 1.0760 ;
      RECT 1.9520 0.8280 2.0020 0.9670 ;
      RECT 1.9520 0.7780 2.0410 0.8280 ;
      RECT 1.9910 0.6280 2.0410 0.7780 ;
      RECT 1.9520 0.5780 2.0410 0.6280 ;
      RECT 1.9520 0.3190 2.0020 0.5780 ;
      RECT 3.8350 0.6670 4.2210 0.7170 ;
      RECT 2.1030 0.6130 2.5490 0.6630 ;
      RECT 2.4330 0.4630 2.4830 0.6130 ;
      RECT 2.4330 0.4130 2.8370 0.4630 ;
      RECT 2.7870 0.4630 2.8370 0.6800 ;
      RECT 2.1030 0.6630 2.1530 0.9120 ;
      RECT 2.1030 0.4130 2.1530 0.6130 ;
      RECT 2.5590 0.7130 2.6850 0.7630 ;
      RECT 2.5590 0.7630 2.6090 0.8670 ;
      RECT 2.6350 0.5630 2.6850 0.7130 ;
      RECT 2.5590 0.8670 2.8530 0.9170 ;
      RECT 2.5430 0.5130 2.6850 0.5630 ;
      RECT 7.6350 1.2000 8.7810 1.2500 ;
      RECT 5.3550 0.6130 6.2570 0.6630 ;
      RECT 6.2070 0.3830 6.2570 0.6130 ;
      RECT 5.5590 0.6630 5.6090 0.9670 ;
      RECT 5.5590 0.9670 6.2570 1.0170 ;
      RECT 6.2070 1.0170 6.2570 1.2400 ;
      RECT 1.6870 0.6780 1.9410 0.7020 ;
      RECT 1.6500 0.7020 1.9410 0.7280 ;
      RECT 1.0230 0.4100 1.3930 0.4600 ;
      RECT 1.3430 0.4600 1.3930 0.5020 ;
      RECT 1.3430 0.5020 1.7370 0.5520 ;
      RECT 1.6870 0.5520 1.7370 0.6780 ;
      RECT 1.6500 0.7280 1.7370 0.7520 ;
      RECT 1.6500 0.7520 1.7000 1.0200 ;
      RECT 1.0230 1.0200 1.7000 1.0700 ;
      RECT 0.8870 0.3100 1.5450 0.3600 ;
      RECT 1.4950 0.3600 1.5450 0.3920 ;
      RECT 0.8870 0.3600 0.9370 0.3920 ;
      RECT 3.7350 0.8670 4.0170 0.9170 ;
      RECT 3.9670 0.9170 4.0170 1.1270 ;
      RECT 3.0150 1.1270 4.0170 1.1770 ;
      RECT 3.0150 1.1770 3.0650 1.2400 ;
      RECT 3.0150 1.0660 3.1150 1.1270 ;
      RECT 3.0650 0.9170 3.1150 1.0660 ;
      RECT 3.0150 0.4130 3.0650 0.8670 ;
      RECT 3.0150 0.8670 3.3090 0.9170 ;
      RECT 3.7350 0.6070 3.7850 0.8670 ;
      RECT 3.7350 0.5570 3.8250 0.6070 ;
      RECT 3.7750 0.4130 3.8250 0.5570 ;
      RECT 1.1750 1.1330 1.5610 1.1830 ;
      RECT 4.4430 0.6130 4.6770 0.6630 ;
      RECT 2.4670 1.5240 4.6770 1.5740 ;
      RECT 2.6190 0.0940 4.3730 0.1440 ;
      RECT 4.2910 0.8670 4.5450 0.9170 ;
      RECT 0.7190 0.5100 1.2570 0.5600 ;
      RECT 6.4190 0.6130 6.7920 0.6630 ;
      RECT 6.7420 0.5700 6.7920 0.6130 ;
      RECT 6.7420 0.5200 7.2270 0.5700 ;
      RECT 7.1770 0.5700 7.2270 0.6040 ;
      RECT 7.1770 0.6040 7.4130 0.6540 ;
      RECT 1.4520 0.6020 1.6370 0.6520 ;
      RECT 0.2050 0.5260 0.2550 0.8410 ;
      RECT 0.2790 0.8910 0.3290 1.2140 ;
      RECT 0.2050 0.4760 0.3290 0.5260 ;
      RECT 0.2790 0.3160 0.3290 0.4760 ;
      RECT 0.2050 0.8410 1.5020 0.8910 ;
      RECT 1.4520 0.6520 1.5020 0.8410 ;
      RECT 8.1830 1.0620 8.6290 1.1120 ;
      RECT 8.1830 0.1260 8.2330 1.0620 ;
      RECT 4.4230 0.0920 6.5020 0.1420 ;
      RECT 4.4230 0.1420 4.4730 0.1940 ;
      RECT 4.3830 0.1940 4.4730 0.2440 ;
      RECT 4.3830 0.2440 4.4330 0.5130 ;
      RECT 4.2310 0.5130 4.4330 0.5630 ;
      RECT 4.2310 0.2770 4.2810 0.5130 ;
      RECT 4.2710 0.5630 4.3210 0.7670 ;
      RECT 4.1910 0.7670 4.3210 0.8170 ;
      RECT 4.1910 0.8170 4.2410 0.9670 ;
      RECT 4.1910 0.9670 4.2810 1.0170 ;
      RECT 4.2310 1.0170 4.2810 1.1900 ;
      RECT 4.2310 1.1900 4.4330 1.2400 ;
      RECT 4.3830 0.9740 4.4330 1.1900 ;
      RECT 0.7190 0.9410 0.9530 0.9910 ;
      RECT 9.2470 0.5890 9.4400 0.6390 ;
      RECT 9.3900 0.5120 9.4400 0.5890 ;
      RECT 9.3900 0.4620 9.5410 0.5120 ;
      RECT 9.3900 0.4120 9.4400 0.4620 ;
      RECT 9.2470 0.3620 9.4400 0.4120 ;
      RECT 9.2470 0.6390 9.2970 0.7720 ;
    LAYER PO ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 3.5570 0.0660 3.5870 0.6370 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 2.7970 0.0660 2.8270 0.6910 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 10.3970 0.0660 10.4270 1.6060 ;
      RECT 4.0130 0.9390 4.0430 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 10.2450 0.0660 10.2750 1.6060 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 5.3810 0.0660 5.4110 0.6910 ;
      RECT 10.0930 0.0660 10.1230 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 9.7890 0.0660 9.8190 1.6060 ;
      RECT 5.8370 0.0660 5.8670 0.7910 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 9.9410 0.0660 9.9710 1.6060 ;
      RECT 9.4850 0.0660 9.5150 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 4.4690 0.0660 4.4990 0.6910 ;
      RECT 4.0130 0.0660 4.0430 0.6370 ;
      RECT 2.7970 0.8390 2.8270 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 5.8370 0.9390 5.8670 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 3.7090 0.0660 3.7390 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 4.4690 0.8390 4.4990 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 9.3330 0.0660 9.3630 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 9.6370 0.0660 9.6670 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 5.3810 0.9590 5.4110 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 7.6610 0.0670 7.6910 1.6050 ;
      RECT 3.5570 0.9390 3.5870 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
    LAYER NWELL ;
      RECT -0.1160 1.5430 10.5730 1.7730 ;
      RECT -0.1160 0.6790 7.5550 1.5430 ;
      RECT 10.3230 0.6790 10.5730 1.5430 ;
      RECT 8.0170 0.4910 9.8630 1.0830 ;
  END
END RSDFFX2_LVT

MACRO SDFFARX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.472 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8390 0.8040 5.2580 0.8540 ;
        RECT 5.1130 0.8540 5.2580 0.9670 ;
        RECT 4.8390 0.8540 4.8890 1.5460 ;
        RECT 5.2080 0.3590 5.2580 0.8040 ;
        RECT 4.8390 0.3090 5.2580 0.3590 ;
        RECT 4.8390 0.1480 4.8890 0.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2650 1.1610 5.3760 1.2210 ;
        RECT 5.1430 1.2210 5.3760 1.2710 ;
        RECT 5.3250 0.2040 5.3750 1.1610 ;
        RECT 5.1430 1.2710 5.1930 1.5460 ;
        RECT 5.1270 0.1540 5.3750 0.2040 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 5.4720 0.0300 ;
        RECT 1.8020 0.0300 1.8520 0.1960 ;
        RECT 1.6470 0.0300 1.6970 0.4080 ;
        RECT 0.5830 0.0300 0.6330 0.5150 ;
        RECT 0.4310 0.0300 0.4810 0.4370 ;
        RECT 4.9910 0.0300 5.0410 0.2330 ;
        RECT 2.7570 0.0300 2.8070 0.2870 ;
        RECT 4.6870 0.0300 4.7370 0.3300 ;
        RECT 1.8020 0.1960 2.1530 0.2460 ;
        RECT 2.7570 0.2870 3.2170 0.3370 ;
        RECT 4.2150 0.3300 4.7530 0.3800 ;
        RECT 2.1030 0.2460 2.1530 0.4500 ;
        RECT 1.9510 0.2460 2.0010 0.4500 ;
        RECT 3.1670 0.3370 3.2170 0.4610 ;
        RECT 3.1670 0.2490 3.2170 0.2870 ;
        RECT 3.1670 0.1990 3.3920 0.2490 ;
    END
  END VSS

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6800 0.7250 0.7300 ;
        RECT 0.4010 0.5530 0.5110 0.6800 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2360 1.3150 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 0.6640 1.0110 0.8150 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 5.4720 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 4.9910 1.0960 5.0410 1.6420 ;
        RECT 1.6470 1.1340 1.6970 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 4.7270 1.3580 4.7770 1.6420 ;
        RECT 3.3430 1.3280 3.3930 1.6420 ;
        RECT 2.1030 1.3640 2.1530 1.6420 ;
        RECT 4.0500 1.3080 4.7770 1.3580 ;
        RECT 3.1500 1.2780 3.3930 1.3280 ;
        RECT 1.9510 1.3140 2.1530 1.3640 ;
        RECT 1.9510 1.0980 2.0010 1.3140 ;
        RECT 2.1030 1.1110 2.1530 1.3140 ;
    END
  END VDD

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9390 0.0880 4.0690 0.1380 ;
        RECT 3.9870 0.1380 4.0690 0.1640 ;
        RECT 2.9390 0.1380 3.0950 0.2070 ;
    END
    ANTENNAGATEAREA 0.0441 ;
  END RSTB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7690 1.4240 1.9410 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  OBS
    LAYER PO ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 2.4930 0.0680 2.5230 0.5420 ;
      RECT 2.4930 0.9900 2.5230 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 4.6210 1.0120 4.6510 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 3.1010 0.0680 3.1310 0.6180 ;
      RECT 4.6210 0.0680 4.6510 0.7870 ;
      RECT 3.7090 0.8820 3.7390 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 5.3810 0.0680 5.4110 1.6060 ;
      RECT 5.2290 0.0680 5.2590 1.6060 ;
      RECT 5.0770 0.0680 5.1070 1.6060 ;
      RECT 4.9250 0.0680 4.9550 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 3.7090 0.0680 3.7390 0.6320 ;
      RECT 4.4690 0.0680 4.4990 1.6060 ;
      RECT 3.1010 0.7580 3.1310 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 4.7730 0.0680 4.8030 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 4.3170 0.0680 4.3470 1.6060 ;
    LAYER NWELL ;
      RECT -0.1150 0.6790 5.5870 1.7730 ;
    LAYER M1 ;
      RECT 1.4520 0.6040 1.6370 0.6540 ;
      RECT 0.2050 0.5280 0.2550 0.8880 ;
      RECT 0.2790 0.9380 0.3290 1.2160 ;
      RECT 0.2050 0.4780 0.3290 0.5280 ;
      RECT 0.2790 0.3180 0.3290 0.4780 ;
      RECT 0.2050 0.8880 1.5020 0.9380 ;
      RECT 1.4520 0.6540 1.5020 0.8880 ;
      RECT 3.4710 1.3080 3.6730 1.3580 ;
      RECT 3.4710 1.1010 3.5210 1.3080 ;
      RECT 3.6230 1.0510 3.6730 1.3080 ;
      RECT 2.7660 1.0010 3.7130 1.0510 ;
      RECT 3.6630 0.5590 3.7130 1.0010 ;
      RECT 3.6230 0.5090 3.7130 0.5590 ;
      RECT 3.6230 0.4700 3.6730 0.5090 ;
      RECT 3.4400 0.4200 3.6730 0.4700 ;
      RECT 3.6230 0.3710 3.6730 0.4200 ;
      RECT 0.7190 0.5120 1.2570 0.5620 ;
      RECT 0.8870 0.3120 1.5450 0.3620 ;
      RECT 0.8870 0.3620 0.9370 0.3940 ;
      RECT 1.4950 0.3620 1.5450 0.3940 ;
      RECT 1.9970 0.0960 2.7070 0.1460 ;
      RECT 4.2710 0.6040 4.9810 0.6540 ;
      RECT 4.2710 0.6540 4.3210 0.9780 ;
      RECT 3.9100 0.9780 4.3210 1.0280 ;
      RECT 3.9100 0.5880 3.9600 0.9780 ;
      RECT 3.9100 0.5380 4.0170 0.5880 ;
      RECT 2.6350 1.4780 3.1570 1.5280 ;
      RECT 2.6350 1.5280 2.6850 1.5650 ;
      RECT 0.7350 1.0420 0.9370 1.0920 ;
      RECT 0.8870 1.0920 0.9370 1.2160 ;
      RECT 0.7350 1.0920 0.7850 1.2160 ;
      RECT 2.3030 1.5260 2.5330 1.5760 ;
      RECT 2.4830 1.4280 2.5330 1.5260 ;
      RECT 2.4830 1.3780 3.2930 1.4280 ;
      RECT 3.2430 1.4280 3.2930 1.5840 ;
      RECT 1.7990 0.6180 2.2450 0.6680 ;
      RECT 1.7990 0.6680 1.8490 0.9140 ;
      RECT 1.7990 0.4220 1.8490 0.6180 ;
      RECT 2.2550 0.5180 2.3810 0.5680 ;
      RECT 2.2550 0.3940 2.3050 0.5180 ;
      RECT 2.3310 0.5680 2.3810 0.7180 ;
      RECT 2.2550 0.7180 2.3810 0.7680 ;
      RECT 2.2550 0.7680 2.3050 0.9140 ;
      RECT 4.2900 1.4290 4.6770 1.4790 ;
      RECT 4.4540 0.7090 4.6770 0.7590 ;
      RECT 4.4540 0.7590 4.5040 1.0990 ;
      RECT 3.8990 1.0990 4.5040 1.1490 ;
      RECT 3.8990 1.1490 3.9490 1.2720 ;
      RECT 3.7230 1.2720 3.9490 1.3220 ;
      RECT 3.7230 1.3220 3.7730 1.5280 ;
      RECT 3.5310 1.5280 3.7730 1.5780 ;
      RECT 1.1750 1.0880 1.5610 1.1380 ;
      RECT 2.6950 1.2780 3.0810 1.3280 ;
      RECT 3.0750 0.7860 3.5970 0.8360 ;
      RECT 3.5470 0.6210 3.5970 0.7860 ;
      RECT 4.3070 0.0880 4.3570 0.2300 ;
      RECT 3.4650 0.2300 4.3570 0.2800 ;
      RECT 3.4650 0.2800 3.5150 0.3140 ;
      RECT 3.3140 0.3140 3.5150 0.3640 ;
      RECT 3.3140 0.3640 3.3640 0.5400 ;
      RECT 3.0750 0.5400 3.3640 0.5900 ;
      RECT 3.6830 0.1880 3.7650 0.2300 ;
      RECT 2.5590 0.6400 3.4610 0.6900 ;
      RECT 2.5590 0.6900 2.6090 1.1580 ;
      RECT 2.5590 0.4840 2.6090 0.6400 ;
      RECT 2.5590 1.2080 2.6090 1.3140 ;
      RECT 2.5590 0.3550 2.6090 0.4340 ;
      RECT 2.5590 1.1580 2.9290 1.2080 ;
      RECT 2.5590 0.4340 2.7770 0.4840 ;
      RECT 2.4070 0.2990 2.4970 0.3810 ;
      RECT 2.4310 0.3810 2.4810 0.9880 ;
      RECT 1.0230 0.9880 2.4810 1.0380 ;
      RECT 2.4070 1.0380 2.4570 1.3140 ;
      RECT 1.3430 0.4620 1.3930 0.5040 ;
      RECT 1.0230 0.4120 1.3930 0.4620 ;
      RECT 1.6500 0.7760 1.7000 0.9880 ;
      RECT 1.6500 0.7260 1.7370 0.7760 ;
      RECT 1.6870 0.5540 1.7370 0.7260 ;
      RECT 1.3430 0.5040 1.7370 0.5540 ;
      RECT 5.0480 0.6040 5.1330 0.6540 ;
      RECT 5.0480 0.5530 5.0980 0.6040 ;
      RECT 5.0480 0.6540 5.0980 0.7040 ;
      RECT 4.4210 0.5030 5.0980 0.5530 ;
      RECT 4.7270 0.7040 5.0980 0.7540 ;
      RECT 4.4210 0.4880 4.4710 0.5030 ;
      RECT 4.7270 0.7540 4.7770 1.2080 ;
      RECT 3.7750 0.4380 4.4710 0.4880 ;
      RECT 4.3670 1.2080 4.7770 1.2580 ;
      RECT 3.7750 0.4880 3.8250 1.1650 ;
      RECT 4.0780 0.4880 4.1280 0.7660 ;
      RECT 4.0780 0.7660 4.2210 0.8160 ;
  END
END SDFFARX1_LVT

MACRO SDFFARX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.776 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.5690 0.0970 5.6790 0.2070 ;
        RECT 5.6110 0.2070 5.6610 0.2700 ;
        RECT 5.2950 0.2700 5.6610 0.3200 ;
        RECT 5.2950 0.1480 5.3450 0.2700 ;
        RECT 5.6110 0.3200 5.6610 0.9180 ;
        RECT 5.2950 0.9180 5.6610 0.9680 ;
        RECT 5.2950 0.9680 5.3450 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 5.7760 0.0300 ;
        RECT 1.8020 0.0300 1.8520 0.1960 ;
        RECT 1.6470 0.0300 1.6970 0.4080 ;
        RECT 0.5830 0.0300 0.6330 0.5150 ;
        RECT 0.4310 0.0300 0.4810 0.4370 ;
        RECT 5.4470 0.0300 5.4970 0.2200 ;
        RECT 4.8390 0.0300 4.8890 0.4080 ;
        RECT 5.1430 0.0300 5.1930 0.3190 ;
        RECT 2.7570 0.0300 2.8070 0.2870 ;
        RECT 4.6870 0.0300 4.7370 0.3300 ;
        RECT 1.8020 0.1960 2.1530 0.2460 ;
        RECT 2.7570 0.2870 3.2170 0.3370 ;
        RECT 4.2150 0.3300 4.7530 0.3800 ;
        RECT 2.1030 0.2460 2.1530 0.4500 ;
        RECT 1.9510 0.2460 2.0010 0.4500 ;
        RECT 3.1670 0.3370 3.2170 0.4610 ;
        RECT 3.1670 0.2490 3.2170 0.2870 ;
        RECT 3.1670 0.1990 3.3920 0.2490 ;
    END
  END VSS

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.9910 0.8040 5.5370 0.8540 ;
        RECT 4.9910 0.8540 5.0410 1.5460 ;
        RECT 5.4870 0.5110 5.5370 0.8040 ;
        RECT 5.4170 0.4440 5.5370 0.5110 ;
        RECT 4.9910 0.3940 5.5370 0.4440 ;
        RECT 4.9910 0.1480 5.0410 0.3940 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6800 0.7250 0.7300 ;
        RECT 0.4010 0.5530 0.5110 0.6800 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2360 1.3150 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 0.6640 1.0110 0.8150 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 5.7760 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 5.4470 1.0520 5.4970 1.6420 ;
        RECT 4.8390 0.9120 4.8890 1.6420 ;
        RECT 5.1430 0.9600 5.1930 1.6420 ;
        RECT 1.6470 1.1340 1.6970 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 4.7270 1.3580 4.7770 1.6420 ;
        RECT 3.3430 1.3280 3.3930 1.6420 ;
        RECT 2.1030 1.3640 2.1530 1.6420 ;
        RECT 4.0500 1.3080 4.7770 1.3580 ;
        RECT 3.1500 1.2780 3.3930 1.3280 ;
        RECT 1.9510 1.3140 2.1530 1.3640 ;
        RECT 1.9510 1.0980 2.0010 1.3140 ;
        RECT 2.1030 1.1110 2.1530 1.3140 ;
    END
  END VDD

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9390 0.0880 4.0690 0.1380 ;
        RECT 3.9870 0.1380 4.0690 0.1740 ;
        RECT 2.9390 0.1380 3.0950 0.2070 ;
    END
    ANTENNAGATEAREA 0.0441 ;
  END RSTB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7690 1.4240 1.9410 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  OBS
    LAYER PO ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 3.7090 0.0680 3.7390 0.6320 ;
      RECT 4.4690 0.0680 4.4990 1.6060 ;
      RECT 3.1010 0.7580 3.1310 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 4.7730 0.0680 4.8030 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 4.3170 0.0680 4.3470 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 2.4930 0.0680 2.5230 0.5420 ;
      RECT 2.4930 0.9900 2.5230 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 4.6210 1.0120 4.6510 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 3.1010 0.0680 3.1310 0.6180 ;
      RECT 4.6210 0.0680 4.6510 0.7870 ;
      RECT 3.7090 0.8820 3.7390 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 5.5330 0.0680 5.5630 1.6060 ;
      RECT 5.3810 0.0680 5.4110 1.6060 ;
      RECT 5.6850 0.0680 5.7150 1.6060 ;
      RECT 5.2290 0.0680 5.2590 1.6060 ;
      RECT 5.0770 0.0680 5.1070 1.6060 ;
      RECT 4.9250 0.0680 4.9550 1.6060 ;
    LAYER NWELL ;
      RECT -0.1150 0.6790 5.8910 1.7730 ;
    LAYER M1 ;
      RECT 5.2000 0.6040 5.4370 0.6540 ;
      RECT 4.7270 0.7540 4.7770 1.2080 ;
      RECT 4.3670 1.2080 4.7770 1.2580 ;
      RECT 4.4210 0.4880 4.4710 0.5030 ;
      RECT 3.7750 0.4380 4.4710 0.4880 ;
      RECT 3.7750 0.4880 3.8250 1.1650 ;
      RECT 4.0780 0.4880 4.1280 0.7660 ;
      RECT 4.0780 0.7660 4.2210 0.8160 ;
      RECT 5.2000 0.6540 5.2500 0.7040 ;
      RECT 5.2000 0.5530 5.2500 0.6040 ;
      RECT 4.4210 0.5030 5.2500 0.5530 ;
      RECT 4.7270 0.7040 5.2500 0.7540 ;
      RECT 1.4520 0.6040 1.6370 0.6540 ;
      RECT 0.2050 0.5280 0.2550 0.8880 ;
      RECT 0.2790 0.9380 0.3290 1.2160 ;
      RECT 0.2050 0.4780 0.3290 0.5280 ;
      RECT 0.2790 0.3180 0.3290 0.4780 ;
      RECT 0.2050 0.8880 1.5020 0.9380 ;
      RECT 1.4520 0.6540 1.5020 0.8880 ;
      RECT 4.4540 0.7090 4.6770 0.7590 ;
      RECT 4.4540 0.7590 4.5040 1.0990 ;
      RECT 3.8990 1.0990 4.5040 1.1490 ;
      RECT 3.8990 1.1490 3.9490 1.2720 ;
      RECT 3.7230 1.2720 3.9490 1.3220 ;
      RECT 3.7230 1.3220 3.7730 1.5280 ;
      RECT 3.5310 1.5280 3.7730 1.5780 ;
      RECT 2.6950 1.2780 3.0810 1.3280 ;
      RECT 3.4710 1.3080 3.6730 1.3580 ;
      RECT 3.4710 1.1010 3.5210 1.3080 ;
      RECT 3.6230 1.0510 3.6730 1.3080 ;
      RECT 2.7660 1.0010 3.7130 1.0510 ;
      RECT 3.6630 0.5590 3.7130 1.0010 ;
      RECT 3.6230 0.5090 3.7130 0.5590 ;
      RECT 3.6230 0.4700 3.6730 0.5090 ;
      RECT 3.4400 0.4200 3.6730 0.4700 ;
      RECT 3.6230 0.3710 3.6730 0.4200 ;
      RECT 0.7190 0.5120 1.2570 0.5620 ;
      RECT 0.8870 0.3120 1.5450 0.3620 ;
      RECT 0.8870 0.3620 0.9370 0.3940 ;
      RECT 1.4950 0.3620 1.5450 0.3940 ;
      RECT 1.9970 0.0960 2.7070 0.1460 ;
      RECT 4.2710 0.6040 5.1330 0.6540 ;
      RECT 4.2710 0.6540 4.3210 0.9780 ;
      RECT 3.9100 0.9780 4.3210 1.0280 ;
      RECT 3.9100 0.5880 3.9600 0.9780 ;
      RECT 3.9100 0.5380 4.0170 0.5880 ;
      RECT 2.6350 1.4780 3.1570 1.5280 ;
      RECT 2.6350 1.5280 2.6850 1.5650 ;
      RECT 0.7350 1.0420 0.9370 1.0920 ;
      RECT 0.8870 1.0920 0.9370 1.2160 ;
      RECT 0.7350 1.0920 0.7850 1.2160 ;
      RECT 2.3030 1.5260 2.5330 1.5760 ;
      RECT 2.4830 1.4280 2.5330 1.5260 ;
      RECT 2.4830 1.3780 3.2930 1.4280 ;
      RECT 3.2430 1.4280 3.2930 1.5840 ;
      RECT 1.7990 0.6180 2.2450 0.6680 ;
      RECT 1.7990 0.6680 1.8490 0.9140 ;
      RECT 1.7990 0.4220 1.8490 0.6180 ;
      RECT 2.2550 0.5180 2.3810 0.5680 ;
      RECT 2.2550 0.3940 2.3050 0.5180 ;
      RECT 2.3310 0.5680 2.3810 0.7180 ;
      RECT 2.2550 0.7180 2.3810 0.7680 ;
      RECT 2.2550 0.7680 2.3050 0.9140 ;
      RECT 4.2900 1.4290 4.6770 1.4790 ;
      RECT 1.1750 1.0880 1.5610 1.1380 ;
      RECT 3.0750 0.7860 3.5970 0.8360 ;
      RECT 3.5470 0.6210 3.5970 0.7860 ;
      RECT 4.3070 0.0880 4.3570 0.2300 ;
      RECT 3.4650 0.2300 4.3570 0.2800 ;
      RECT 3.6830 0.2800 3.7650 0.2900 ;
      RECT 3.4650 0.2800 3.5150 0.3140 ;
      RECT 3.3140 0.3140 3.5150 0.3640 ;
      RECT 3.3140 0.3640 3.3640 0.5400 ;
      RECT 3.0750 0.5400 3.3640 0.5900 ;
      RECT 3.6830 0.1880 3.7650 0.2300 ;
      RECT 2.5590 0.6400 3.4610 0.6900 ;
      RECT 2.5590 0.6900 2.6090 1.1580 ;
      RECT 2.5590 0.4840 2.6090 0.6400 ;
      RECT 2.5590 1.2080 2.6090 1.3140 ;
      RECT 2.5590 0.3550 2.6090 0.4340 ;
      RECT 2.5590 1.1580 2.9290 1.2080 ;
      RECT 2.5590 0.4340 2.7770 0.4840 ;
      RECT 2.4070 0.2990 2.4970 0.3810 ;
      RECT 2.4310 0.3810 2.4810 0.9880 ;
      RECT 1.0230 0.9880 2.4810 1.0380 ;
      RECT 2.4070 1.0380 2.4570 1.3140 ;
      RECT 1.3430 0.4620 1.3930 0.5040 ;
      RECT 1.0230 0.4120 1.3930 0.4620 ;
      RECT 1.6500 0.7760 1.7000 0.9880 ;
      RECT 1.6500 0.7260 1.7370 0.7760 ;
      RECT 1.6870 0.5540 1.7370 0.7260 ;
      RECT 1.3430 0.5040 1.7370 0.5540 ;
  END
END SDFFARX2_LVT

MACRO SDFFASRSX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.08 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.7510 1.2210 6.0250 1.2710 ;
        RECT 5.7510 1.2710 5.8010 1.5460 ;
        RECT 5.8730 1.1610 6.0250 1.2210 ;
        RECT 5.9750 0.2040 6.0250 1.1610 ;
        RECT 5.7350 0.1540 6.0250 0.2040 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 6.0800 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 1.6470 1.1340 1.6970 1.6420 ;
        RECT 5.2950 0.9470 5.3450 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 5.5990 1.1860 5.6490 1.6420 ;
        RECT 5.0310 1.3580 5.0810 1.6420 ;
        RECT 3.3430 1.3280 3.3930 1.6420 ;
        RECT 2.1030 1.3540 2.1530 1.6420 ;
        RECT 4.2020 1.3080 5.0810 1.3580 ;
        RECT 3.1500 1.2780 3.5520 1.3280 ;
        RECT 1.9510 1.3040 2.1530 1.3540 ;
        RECT 1.9510 1.0880 2.0010 1.3040 ;
        RECT 2.1030 1.1010 2.1530 1.3040 ;
    END
  END VDD

  PIN SO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.1430 0.8220 5.8250 0.8720 ;
        RECT 5.5690 0.8720 5.6790 0.9670 ;
        RECT 5.1430 0.8720 5.1930 1.5460 ;
        RECT 5.7750 0.4300 5.8250 0.8220 ;
        RECT 5.1430 0.3800 5.8250 0.4300 ;
        RECT 5.1430 0.1480 5.1930 0.3800 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END SO

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 0.6640 1.0110 0.8150 ;
    END
    ANTENNAGATEAREA 0.0255 ;
  END D

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9390 0.0880 4.2210 0.1380 ;
        RECT 4.1390 0.1380 4.2210 0.1640 ;
        RECT 2.9390 0.1380 3.0950 0.2070 ;
    END
    ANTENNAGATEAREA 0.039 ;
  END RSTB

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6800 0.7250 0.7300 ;
        RECT 0.4010 0.5530 0.5110 0.6800 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2360 1.3150 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.7470 0.8190 4.9190 0.9960 ;
    END
    ANTENNAGATEAREA 0.039 ;
  END SETB

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 6.0800 0.0300 ;
        RECT 1.6470 0.0300 1.6970 0.1960 ;
        RECT 5.2950 0.0300 5.3450 0.2200 ;
        RECT 0.5830 0.0300 0.6330 0.5150 ;
        RECT 0.4310 0.0300 0.4810 0.4370 ;
        RECT 5.5990 0.0300 5.6490 0.2200 ;
        RECT 2.7570 0.0300 2.8070 0.2870 ;
        RECT 4.9910 0.0300 5.0410 0.3300 ;
        RECT 1.6470 0.1960 2.1530 0.2460 ;
        RECT 2.7570 0.2870 3.3690 0.3370 ;
        RECT 4.3670 0.3300 5.0570 0.3800 ;
        RECT 2.1030 0.2460 2.1530 0.4500 ;
        RECT 1.9510 0.2460 2.0010 0.4500 ;
        RECT 1.6470 0.2460 1.6970 0.4080 ;
        RECT 3.3190 0.3370 3.3690 0.4610 ;
        RECT 3.1670 0.3370 3.2170 0.4610 ;
    END
  END VSS

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7690 1.4240 1.9410 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4470 1.0590 5.8310 1.0670 ;
        RECT 5.7210 1.0670 5.8310 1.1190 ;
        RECT 5.4470 1.0170 5.9250 1.0590 ;
        RECT 5.4470 1.0670 5.4970 1.5460 ;
        RECT 5.7210 1.0090 5.9250 1.0170 ;
        RECT 5.8750 0.3200 5.9250 1.0090 ;
        RECT 5.4470 0.2700 5.9250 0.3200 ;
        RECT 5.4470 0.1480 5.4970 0.2700 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q
  OBS
    LAYER PO ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 3.1010 0.7580 3.1310 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 5.3810 0.0680 5.4110 1.6060 ;
      RECT 5.8370 0.0680 5.8670 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 4.3170 0.0680 4.3470 1.6060 ;
      RECT 4.7730 0.0680 4.8030 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 3.7090 0.0680 3.7390 1.6060 ;
      RECT 4.4690 0.0680 4.4990 1.6060 ;
      RECT 5.6850 0.0680 5.7150 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 4.6210 0.0680 4.6510 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 5.5330 0.0680 5.5630 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 5.0770 0.0680 5.1070 1.6060 ;
      RECT 2.4930 0.0680 2.5230 0.5420 ;
      RECT 5.9890 0.0680 6.0190 1.6060 ;
      RECT 2.4930 0.9900 2.5230 1.6060 ;
      RECT 4.9250 0.0680 4.9550 0.7870 ;
      RECT 3.1010 0.0680 3.1310 0.6180 ;
      RECT 3.8610 0.8820 3.8910 1.6060 ;
      RECT 5.2290 0.0680 5.2590 1.6060 ;
      RECT 4.9250 0.9120 4.9550 1.6060 ;
      RECT 3.8610 0.0680 3.8910 0.6320 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
    LAYER NWELL ;
      RECT -0.1150 0.6790 6.1950 1.7730 ;
    LAYER M1 ;
      RECT 2.7660 0.9560 3.8650 1.0060 ;
      RECT 3.7750 1.0060 3.8650 1.0510 ;
      RECT 3.8150 0.6560 3.8650 0.9560 ;
      RECT 3.7750 1.0510 3.8250 1.3080 ;
      RECT 3.7750 0.6060 3.8650 0.6560 ;
      RECT 3.6230 1.3080 3.8250 1.3580 ;
      RECT 3.7750 0.4960 3.8250 0.6060 ;
      RECT 3.6230 1.2160 3.6730 1.3080 ;
      RECT 3.6230 0.4460 3.8250 0.4960 ;
      RECT 3.3020 1.1660 3.6730 1.2160 ;
      RECT 3.6230 0.3710 3.6730 0.4460 ;
      RECT 3.7750 0.3710 3.8250 0.4460 ;
      RECT 2.5590 0.6400 3.4610 0.6900 ;
      RECT 2.5590 0.6900 2.6090 1.1580 ;
      RECT 2.5590 0.4840 2.6090 0.6400 ;
      RECT 2.5590 1.2080 2.6090 1.3140 ;
      RECT 2.5590 0.3550 2.6090 0.4340 ;
      RECT 2.5590 1.1580 2.9290 1.2080 ;
      RECT 2.5590 0.4340 2.7770 0.4840 ;
      RECT 2.4070 0.2990 2.4970 0.3810 ;
      RECT 2.4310 0.3810 2.4810 0.9880 ;
      RECT 2.4070 1.0380 2.4570 1.3140 ;
      RECT 1.0230 0.9880 2.4810 1.0380 ;
      RECT 1.3430 0.4620 1.3930 0.5040 ;
      RECT 1.0230 0.4120 1.3930 0.4620 ;
      RECT 1.6500 0.7760 1.7000 0.9880 ;
      RECT 1.6500 0.7260 1.7370 0.7760 ;
      RECT 1.6870 0.5540 1.7370 0.7260 ;
      RECT 1.3430 0.5040 1.7370 0.5540 ;
      RECT 3.0750 0.7860 3.7650 0.8360 ;
      RECT 2.3150 1.5260 2.5330 1.5760 ;
      RECT 2.4830 1.4280 2.5330 1.5260 ;
      RECT 2.4830 1.3780 3.2930 1.4280 ;
      RECT 3.2430 1.4280 3.2930 1.5440 ;
      RECT 4.5610 0.7090 4.9810 0.7590 ;
      RECT 4.5610 0.7590 4.6110 1.0990 ;
      RECT 4.0510 1.0990 4.6110 1.1490 ;
      RECT 4.0510 1.1490 4.1010 1.2720 ;
      RECT 3.8750 1.2720 4.1010 1.3220 ;
      RECT 3.8750 1.3220 3.9250 1.4280 ;
      RECT 3.6830 1.4280 3.9250 1.4780 ;
      RECT 4.5190 1.2080 4.9050 1.2580 ;
      RECT 2.6950 1.2780 3.0810 1.3280 ;
      RECT 4.4230 0.6040 5.5890 0.6540 ;
      RECT 4.4230 0.6540 4.4730 0.9780 ;
      RECT 4.0620 0.9780 4.4730 1.0280 ;
      RECT 4.0620 0.4960 4.1120 0.9780 ;
      RECT 4.0620 0.4460 4.1690 0.4960 ;
      RECT 4.4420 1.4080 4.9810 1.4580 ;
      RECT 2.6350 1.4780 3.1570 1.5280 ;
      RECT 2.6350 1.5280 2.6850 1.5650 ;
      RECT 0.8870 0.3120 1.5450 0.3620 ;
      RECT 0.8870 0.3620 0.9370 0.3940 ;
      RECT 1.4950 0.3620 1.5450 0.3940 ;
      RECT 1.7990 0.6180 2.2450 0.6680 ;
      RECT 1.7990 0.6680 1.8490 0.9140 ;
      RECT 1.7990 0.4220 1.8490 0.6180 ;
      RECT 2.2550 0.5180 2.3810 0.5680 ;
      RECT 2.2550 0.3940 2.3050 0.5180 ;
      RECT 2.3310 0.5680 2.3810 0.7180 ;
      RECT 2.2550 0.7180 2.3810 0.7680 ;
      RECT 2.2550 0.7680 2.3050 0.9140 ;
      RECT 0.7350 1.0420 0.9370 1.0920 ;
      RECT 0.8870 1.0920 0.9370 1.2160 ;
      RECT 0.7350 1.0920 0.7850 1.2160 ;
      RECT 0.7190 0.5120 1.2570 0.5620 ;
      RECT 2.0110 0.0960 2.7070 0.1460 ;
      RECT 1.1750 1.0880 1.5610 1.1380 ;
      RECT 3.5020 1.5280 4.8420 1.5780 ;
      RECT 5.0310 0.7040 5.7250 0.7540 ;
      RECT 5.6750 0.5540 5.7250 0.7040 ;
      RECT 4.6780 0.5040 5.7250 0.5540 ;
      RECT 5.0310 0.7540 5.0810 1.1080 ;
      RECT 4.6710 1.1080 5.0810 1.1580 ;
      RECT 4.6780 0.4880 4.7280 0.5040 ;
      RECT 4.2300 0.4380 4.7280 0.4880 ;
      RECT 4.2300 0.7660 4.3730 0.8160 ;
      RECT 4.2300 0.4880 4.2800 0.7660 ;
      RECT 4.2300 0.3960 4.2800 0.4380 ;
      RECT 3.9270 0.3460 4.2800 0.3960 ;
      RECT 3.9270 0.3960 3.9770 1.1650 ;
      RECT 1.4520 0.6040 1.6370 0.6540 ;
      RECT 0.2050 0.5280 0.2550 0.8880 ;
      RECT 0.2790 0.9380 0.3290 1.2160 ;
      RECT 0.2050 0.4780 0.3290 0.5280 ;
      RECT 0.2790 0.3180 0.3290 0.4780 ;
      RECT 0.2050 0.8880 1.5020 0.9380 ;
      RECT 1.4520 0.6540 1.5020 0.8880 ;
      RECT 4.4590 0.0880 4.5090 0.2300 ;
      RECT 3.5110 0.2300 4.5090 0.2800 ;
      RECT 3.5110 0.2800 3.5610 0.5400 ;
      RECT 3.0750 0.5400 3.5610 0.5900 ;
      RECT 3.8350 0.1880 3.9170 0.2300 ;
  END
END SDFFASRSX1_LVT

MACRO RSDFFNSRASRNX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.336 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 10.3360 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 2.1030 1.1310 2.1530 1.6420 ;
        RECT 1.7990 1.1310 1.8490 1.6420 ;
        RECT 1.6470 1.1310 1.6970 1.6420 ;
        RECT 8.3750 1.4540 8.4250 1.6420 ;
        RECT 3.9670 1.2700 4.0170 1.6420 ;
        RECT 2.2550 1.2940 2.3050 1.6420 ;
        RECT 5.7510 1.4040 8.4250 1.4540 ;
        RECT 3.7580 1.2200 5.0570 1.2700 ;
        RECT 2.2550 1.2440 2.7770 1.2940 ;
        RECT 5.7510 1.2790 5.8010 1.4040 ;
        RECT 6.9670 0.9590 7.0170 1.4040 ;
        RECT 6.5110 0.9530 6.5610 1.4040 ;
    END
  END VDD

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.8150 0.4010 7.5150 0.4510 ;
        RECT 6.8150 0.1570 6.8650 0.4010 ;
        RECT 7.3930 0.4510 7.5150 0.5110 ;
        RECT 7.1190 0.1570 7.1690 0.4010 ;
        RECT 7.4650 0.5110 7.5150 0.8590 ;
        RECT 6.8150 0.8590 7.5150 0.9090 ;
        RECT 6.8150 0.9090 6.8650 1.3090 ;
        RECT 7.1190 0.9090 7.1690 1.3090 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END QN

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 10.3360 0.0300 ;
        RECT 2.1030 0.0300 2.1530 0.3070 ;
        RECT 9.3990 0.0300 9.4490 0.4260 ;
        RECT 1.6470 0.0300 1.6970 0.4050 ;
        RECT 6.9670 0.0300 7.0170 0.2410 ;
        RECT 1.7990 0.0300 1.8490 0.4050 ;
        RECT 8.0310 0.0300 8.0810 0.4260 ;
        RECT 0.5830 0.0300 0.6330 0.5120 ;
        RECT 0.4310 0.0300 0.4810 0.4340 ;
        RECT 8.9430 0.0300 8.9930 0.1980 ;
        RECT 6.6870 0.0300 6.7370 0.2880 ;
        RECT 2.1030 0.3070 3.9770 0.3570 ;
        RECT 5.7350 0.2880 6.7370 0.3380 ;
        RECT 2.5590 0.3570 2.6090 0.5570 ;
        RECT 3.7750 0.3570 3.8250 0.5570 ;
        RECT 2.7110 0.3570 2.7610 0.5570 ;
        RECT 3.9270 0.3570 3.9770 0.5330 ;
        RECT 2.1030 0.3570 2.1530 0.4050 ;
        RECT 3.9270 0.2380 3.9770 0.3070 ;
        RECT 3.9270 0.1880 5.0570 0.2380 ;
        RECT 4.3830 0.2380 4.4330 0.3490 ;
    END
  END VSS

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.9790 0.8570 6.1350 0.9750 ;
        RECT 5.9790 0.9750 6.0290 1.0790 ;
        RECT 5.4470 1.0790 6.0290 1.1290 ;
        RECT 5.4470 1.1290 5.4970 1.3200 ;
        RECT 4.1550 1.3200 5.4970 1.3700 ;
        RECT 4.1550 1.3700 4.2050 1.4550 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.5470 0.0880 6.4850 0.0970 ;
        RECT 3.4390 0.0970 6.4850 0.1380 ;
        RECT 3.4390 0.1380 3.5970 0.2100 ;
        RECT 6.4350 0.1380 6.4850 0.1700 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3770 1.4650 2.5490 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.5210 0.2490 9.6310 0.3590 ;
        RECT 9.5320 0.3590 9.5820 0.5270 ;
        RECT 9.3070 0.5270 9.5820 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6570 0.7050 4.8130 0.7310 ;
        RECT 4.6570 0.7310 5.1170 0.7810 ;
        RECT 4.7630 0.5970 4.8130 0.7050 ;
        RECT 4.6570 0.7810 4.8130 0.8150 ;
        RECT 5.0670 0.7810 5.1170 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 8.0150 0.9420 9.6330 1.0020 ;
        RECT 9.5230 0.6900 9.6330 0.9420 ;
        RECT 9.3990 0.6270 9.4490 0.9420 ;
    END
  END VDDG

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2520 1.3330 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6780 0.7250 0.7280 ;
        RECT 0.4010 0.5510 0.5110 0.6780 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 1.1610 1.0110 1.3160 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D
  OBS
    LAYER M1 ;
      RECT 4.8230 1.1200 5.3450 1.1700 ;
      RECT 4.2130 0.8580 4.3730 0.9080 ;
      RECT 4.2130 0.9080 4.2630 0.9680 ;
      RECT 3.6830 0.9680 4.2630 1.0180 ;
      RECT 1.4520 0.6020 1.6370 0.6520 ;
      RECT 0.2050 0.8410 1.5020 0.8910 ;
      RECT 1.4520 0.6520 1.5020 0.8410 ;
      RECT 0.2050 0.5260 0.2550 0.8410 ;
      RECT 0.2790 0.8910 0.3290 1.2140 ;
      RECT 0.2050 0.4760 0.3290 0.5260 ;
      RECT 0.2790 0.3160 0.3290 0.4760 ;
      RECT 3.1670 0.8540 4.0690 0.9040 ;
      RECT 3.1670 0.6130 3.2170 0.8540 ;
      RECT 3.1670 0.9040 3.2170 1.0590 ;
      RECT 3.1670 0.5630 3.3690 0.6130 ;
      RECT 3.1670 1.0590 3.5370 1.1090 ;
      RECT 3.3190 0.4070 3.3690 0.5630 ;
      RECT 3.1670 0.4130 3.2170 0.5630 ;
      RECT 3.1670 1.1090 3.2170 1.3370 ;
      RECT 6.5870 0.6420 7.1090 0.6920 ;
      RECT 5.9430 0.4500 5.9930 0.7290 ;
      RECT 5.9430 0.7290 6.3090 0.7790 ;
      RECT 6.2590 0.7790 6.3090 1.1790 ;
      RECT 5.5990 0.4000 6.6370 0.4500 ;
      RECT 6.5870 0.4500 6.6370 0.6420 ;
      RECT 5.6000 1.1790 6.3090 1.2290 ;
      RECT 5.5990 0.2970 5.6490 0.4000 ;
      RECT 5.5990 0.4500 5.6490 0.5630 ;
      RECT 5.6000 1.2290 5.6500 1.3530 ;
      RECT 5.1470 0.1880 5.7410 0.2380 ;
      RECT 5.1470 0.2380 5.1970 0.2880 ;
      RECT 4.5060 0.2880 5.1970 0.3380 ;
      RECT 4.1190 0.4550 4.1690 0.6130 ;
      RECT 3.6830 0.6130 4.1690 0.6630 ;
      RECT 4.5060 0.3380 4.5560 0.4050 ;
      RECT 4.1190 0.4050 4.5560 0.4550 ;
      RECT 3.0150 0.8130 3.1050 0.8630 ;
      RECT 3.0550 0.4620 3.1050 0.8130 ;
      RECT 3.0150 0.8630 3.0650 1.0830 ;
      RECT 2.9990 0.4120 3.1050 0.4620 ;
      RECT 2.2550 1.0830 3.0650 1.1330 ;
      RECT 3.0150 1.1330 3.0650 1.3540 ;
      RECT 2.2550 0.7520 2.3050 1.0830 ;
      RECT 2.2550 0.7020 2.3450 0.7520 ;
      RECT 2.2950 0.5510 2.3450 0.7020 ;
      RECT 2.2550 0.5010 2.3450 0.5510 ;
      RECT 2.2550 0.4070 2.3050 0.5010 ;
      RECT 2.4070 0.6130 2.8530 0.6630 ;
      RECT 2.4070 0.6630 2.4570 1.0040 ;
      RECT 2.4070 0.4130 2.4570 0.6130 ;
      RECT 8.3190 0.8200 8.8670 0.8700 ;
      RECT 1.6500 0.7020 1.9410 0.7280 ;
      RECT 1.6870 0.6780 1.9410 0.7020 ;
      RECT 1.3430 0.4600 1.3930 0.5020 ;
      RECT 1.0230 0.4100 1.3930 0.4600 ;
      RECT 1.0230 1.0200 1.7000 1.0700 ;
      RECT 1.6500 0.7520 1.7000 1.0200 ;
      RECT 1.6500 0.7280 1.7370 0.7520 ;
      RECT 1.6870 0.5520 1.7370 0.6780 ;
      RECT 1.3430 0.5020 1.7370 0.5520 ;
      RECT 0.8870 0.3100 1.5450 0.3600 ;
      RECT 1.4950 0.3600 1.5450 0.3920 ;
      RECT 0.8870 0.3600 0.9370 0.3920 ;
      RECT 5.6590 0.8660 5.8080 0.9160 ;
      RECT 5.7580 0.9160 5.8080 0.9670 ;
      RECT 5.7580 0.9670 5.8930 1.0170 ;
      RECT 7.1680 0.6130 7.4130 0.6630 ;
      RECT 6.3590 0.8090 6.4090 1.3010 ;
      RECT 6.3590 0.5500 6.4090 0.7590 ;
      RECT 6.1310 0.5000 6.4090 0.5500 ;
      RECT 6.1310 0.5500 6.1810 0.6790 ;
      RECT 6.6630 0.8090 6.7130 1.3010 ;
      RECT 7.1680 0.6630 7.2180 0.7590 ;
      RECT 6.3590 0.7590 7.2180 0.8090 ;
      RECT 1.9910 0.6280 2.2450 0.6520 ;
      RECT 1.9520 0.6020 2.2450 0.6280 ;
      RECT 1.9910 0.6520 2.0410 0.7780 ;
      RECT 1.9520 0.5780 2.0410 0.6020 ;
      RECT 1.9520 0.7780 2.0410 0.8280 ;
      RECT 1.9520 0.3190 2.0020 0.5780 ;
      RECT 1.9520 0.8280 2.0020 1.0760 ;
      RECT 8.6230 0.7090 9.1610 0.7590 ;
      RECT 4.6710 0.4880 5.2330 0.5380 ;
      RECT 5.1830 0.5380 5.2330 1.0200 ;
      RECT 4.6870 1.0200 5.2330 1.0700 ;
      RECT 4.4230 0.7880 4.4730 1.1200 ;
      RECT 3.3740 0.7380 4.4750 0.7880 ;
      RECT 4.2310 0.5050 4.2810 0.7380 ;
      RECT 4.6870 1.0700 4.7370 1.1200 ;
      RECT 3.9110 1.1200 4.7370 1.1700 ;
      RECT 5.2010 1.5200 8.3250 1.5700 ;
      RECT 9.2470 0.6770 9.2970 0.7680 ;
      RECT 9.2070 0.4270 9.2970 0.4620 ;
      RECT 9.2470 0.1260 9.2970 0.4270 ;
      RECT 9.2070 0.6270 9.2970 0.6770 ;
      RECT 9.2070 0.5120 9.2570 0.6270 ;
      RECT 9.0030 0.4770 9.2570 0.5120 ;
      RECT 9.0030 0.4620 9.2970 0.4770 ;
      RECT 2.9220 0.0940 3.3150 0.1440 ;
      RECT 4.4430 1.5200 5.1330 1.5700 ;
      RECT 4.8980 0.6130 5.1330 0.6630 ;
      RECT 5.4470 0.8670 5.5890 0.9170 ;
      RECT 5.4470 0.6630 5.4970 0.8670 ;
      RECT 5.4470 0.6130 5.8930 0.6630 ;
      RECT 4.5350 0.9200 4.9650 0.9700 ;
      RECT 4.9150 0.8310 4.9650 0.9200 ;
      RECT 4.5350 0.9700 4.5850 1.0340 ;
      RECT 4.5350 0.5050 4.5850 0.9200 ;
      RECT 4.2910 1.4200 5.5970 1.4700 ;
      RECT 3.3030 1.1900 3.6890 1.2400 ;
      RECT 5.8800 1.2870 6.2730 1.3370 ;
      RECT 3.2270 1.3890 3.7650 1.4390 ;
      RECT 2.6190 1.5240 3.9170 1.5740 ;
      RECT 7.3310 1.1990 8.6290 1.2490 ;
      RECT 7.9390 0.5270 8.5370 0.5770 ;
      RECT 8.4870 0.5770 8.5370 0.7700 ;
      RECT 8.4870 0.3480 8.5370 0.5270 ;
      RECT 8.1830 0.5770 8.2330 0.8720 ;
      RECT 8.1830 0.1260 8.2330 0.5270 ;
      RECT 8.6230 0.1320 8.8570 0.1820 ;
      RECT 7.8790 1.0620 8.3280 1.1120 ;
      RECT 7.8790 0.6770 7.9290 1.0620 ;
      RECT 7.8390 0.6270 7.9290 0.6770 ;
      RECT 7.8390 0.4770 7.8890 0.6270 ;
      RECT 7.8390 0.4270 7.9290 0.4770 ;
      RECT 7.8790 0.1260 7.9290 0.4270 ;
      RECT 0.7190 0.5100 1.2570 0.5600 ;
      RECT 1.1750 1.1330 1.5610 1.1830 ;
      RECT 0.7190 0.9410 0.9530 0.9910 ;
      RECT 8.8510 1.0620 9.3890 1.1120 ;
      RECT 8.3190 0.2480 9.1610 0.2980 ;
      RECT 2.8630 0.7130 2.9890 0.7630 ;
      RECT 2.8630 0.7630 2.9130 1.0330 ;
      RECT 2.9390 0.5630 2.9890 0.7130 ;
      RECT 2.8470 0.5130 2.9890 0.5630 ;
      RECT 4.8230 0.3880 5.4970 0.4380 ;
      RECT 5.4470 0.4380 5.4970 0.5630 ;
      RECT 5.4470 0.2970 5.4970 0.3880 ;
      RECT 5.2950 0.9670 5.5130 1.0170 ;
      RECT 5.2950 0.4380 5.3450 0.9670 ;
      RECT 5.2950 1.0170 5.3450 1.1200 ;
      RECT 5.2950 1.1700 5.3450 1.2700 ;
    LAYER PO ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 5.8370 0.0660 5.8670 0.6910 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 3.1010 0.8400 3.1310 1.6060 ;
      RECT 5.8370 0.9390 5.8670 1.6060 ;
      RECT 5.5330 0.0660 5.5630 0.6370 ;
      RECT 3.1010 0.0660 3.1310 0.6370 ;
      RECT 3.7090 0.0660 3.7390 0.6910 ;
      RECT 9.3330 0.0660 9.3630 1.6060 ;
      RECT 5.0770 0.0660 5.1070 0.6910 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 9.6370 0.0660 9.6670 1.6060 ;
      RECT 4.7730 0.8920 4.8030 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 5.5330 0.8390 5.5630 1.6060 ;
      RECT 9.7890 0.0660 9.8190 1.6060 ;
      RECT 10.2450 0.0660 10.2750 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 9.9410 0.0660 9.9710 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 10.0930 0.0660 10.1230 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 4.7730 0.0660 4.8030 0.6910 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 3.7090 0.9390 3.7390 1.6060 ;
      RECT 7.3570 0.0670 7.3870 1.6050 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 5.0770 0.8390 5.1070 1.6060 ;
      RECT 9.4850 0.0660 9.5150 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
    LAYER NWELL ;
      RECT 7.7120 0.4910 9.7230 1.0830 ;
      RECT -0.1150 1.5430 10.4580 1.7730 ;
      RECT -0.1150 0.6790 7.2500 1.5430 ;
      RECT 10.1830 0.6790 10.4580 1.5430 ;
  END
END RSDFFNSRASRNX2_LVT

MACRO RSDFFNSRASRQX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.184 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 10.1840 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 2.1030 1.1310 2.1530 1.6420 ;
        RECT 1.7990 1.1310 1.8490 1.6420 ;
        RECT 1.6470 1.1310 1.6970 1.6420 ;
        RECT 8.2230 1.4540 8.2730 1.6420 ;
        RECT 3.9670 1.2700 4.0170 1.6420 ;
        RECT 2.2550 1.2940 2.3050 1.6420 ;
        RECT 5.7510 1.4040 8.2730 1.4540 ;
        RECT 3.7580 1.2200 5.0570 1.2700 ;
        RECT 2.2550 1.2440 2.7770 1.2940 ;
        RECT 5.7510 1.2790 5.8010 1.4040 ;
        RECT 6.8150 0.9590 6.8650 1.4040 ;
        RECT 6.5110 0.9530 6.5610 1.4040 ;
    END
  END VDD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.9670 0.9690 7.5010 1.0190 ;
        RECT 7.4510 0.3510 7.5010 0.9690 ;
        RECT 6.9670 1.0190 7.1990 1.1290 ;
        RECT 6.9510 0.3010 7.5010 0.3510 ;
        RECT 6.9670 1.1290 7.0170 1.3270 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 10.1840 0.0300 ;
        RECT 2.1030 0.0300 2.1530 0.3070 ;
        RECT 9.2470 0.0300 9.2970 0.4260 ;
        RECT 1.6470 0.0300 1.6970 0.4050 ;
        RECT 6.8150 0.0300 6.8650 0.2410 ;
        RECT 1.7990 0.0300 1.8490 0.4050 ;
        RECT 7.8790 0.0300 7.9290 0.4260 ;
        RECT 0.5830 0.0300 0.6330 0.5120 ;
        RECT 0.4310 0.0300 0.4810 0.4340 ;
        RECT 8.7910 0.0300 8.8410 0.1980 ;
        RECT 6.6870 0.0300 6.7370 0.2880 ;
        RECT 2.1030 0.3070 3.9770 0.3570 ;
        RECT 5.7350 0.2880 6.7370 0.3380 ;
        RECT 2.5590 0.3570 2.6090 0.5570 ;
        RECT 3.7750 0.3570 3.8250 0.5570 ;
        RECT 2.7110 0.3570 2.7610 0.5570 ;
        RECT 3.9270 0.3570 3.9770 0.5330 ;
        RECT 2.1030 0.3570 2.1530 0.4050 ;
        RECT 3.9270 0.2380 3.9770 0.3070 ;
        RECT 3.9270 0.1880 5.0570 0.2380 ;
        RECT 4.3830 0.2380 4.4330 0.3490 ;
    END
  END VSS

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.9790 0.8570 6.1350 0.9750 ;
        RECT 5.9790 0.9750 6.0290 1.0790 ;
        RECT 5.4470 1.0790 6.0290 1.1290 ;
        RECT 5.4470 1.1290 5.4970 1.3200 ;
        RECT 4.1550 1.3200 5.4970 1.3700 ;
        RECT 4.1550 1.3700 4.2050 1.4550 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.5470 0.0880 6.4850 0.0970 ;
        RECT 3.4390 0.0970 6.4850 0.1380 ;
        RECT 3.4390 0.1380 3.5970 0.2100 ;
        RECT 6.4350 0.1380 6.4850 0.1700 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3770 1.4650 2.5490 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.3690 0.2490 9.4790 0.3590 ;
        RECT 9.3800 0.3590 9.4300 0.4960 ;
        RECT 9.1550 0.4960 9.4300 0.5460 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6570 0.7310 5.1170 0.7810 ;
        RECT 4.6570 0.7050 4.8130 0.7310 ;
        RECT 4.6570 0.7810 4.8130 0.8150 ;
        RECT 5.0670 0.7810 5.1170 0.9330 ;
        RECT 4.7630 0.5970 4.8130 0.7050 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 7.8630 0.9420 9.4810 1.0020 ;
        RECT 9.3710 0.6900 9.4810 0.9420 ;
        RECT 9.2470 0.6270 9.2970 0.9420 ;
    END
  END VDDG

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2520 1.3330 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6780 0.7250 0.7280 ;
        RECT 0.4010 0.5510 0.5110 0.6780 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 1.1610 1.0110 1.3160 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D
  OBS
    LAYER M1 ;
      RECT 0.2790 0.3160 0.3290 0.4760 ;
      RECT 3.1670 0.8540 4.0690 0.9040 ;
      RECT 3.1670 0.6130 3.2170 0.8540 ;
      RECT 3.1670 0.9040 3.2170 1.0590 ;
      RECT 3.1670 0.5630 3.3690 0.6130 ;
      RECT 3.1670 1.0590 3.5370 1.1090 ;
      RECT 3.3190 0.4070 3.3690 0.5630 ;
      RECT 3.1670 0.4130 3.2170 0.5630 ;
      RECT 3.1670 1.1090 3.2170 1.3370 ;
      RECT 5.5990 0.4000 6.6370 0.4500 ;
      RECT 6.5870 0.4500 6.6370 0.6920 ;
      RECT 5.9430 0.4500 5.9930 0.7290 ;
      RECT 5.9430 0.7290 6.3090 0.7790 ;
      RECT 6.2590 0.7790 6.3090 1.1790 ;
      RECT 5.6000 1.1790 6.3090 1.2290 ;
      RECT 5.5990 0.4500 5.6490 0.5630 ;
      RECT 5.5990 0.2970 5.6490 0.4000 ;
      RECT 5.6000 1.2290 5.6500 1.3530 ;
      RECT 3.0550 0.4620 3.1050 0.8130 ;
      RECT 2.9990 0.4120 3.1050 0.4620 ;
      RECT 3.0150 0.8130 3.1050 0.8630 ;
      RECT 3.0150 0.8630 3.0650 1.0830 ;
      RECT 2.2550 1.0830 3.0650 1.1330 ;
      RECT 3.0150 1.1330 3.0650 1.3540 ;
      RECT 2.2550 0.7520 2.3050 1.0830 ;
      RECT 2.2550 0.7020 2.3450 0.7520 ;
      RECT 2.2950 0.5510 2.3450 0.7020 ;
      RECT 2.2550 0.5010 2.3450 0.5510 ;
      RECT 2.2550 0.4070 2.3050 0.5010 ;
      RECT 2.4070 0.6130 2.8530 0.6630 ;
      RECT 2.4070 0.6630 2.4570 1.0040 ;
      RECT 2.4070 0.4130 2.4570 0.6130 ;
      RECT 8.1670 0.8200 8.7150 0.8700 ;
      RECT 1.6500 0.7020 1.9410 0.7280 ;
      RECT 1.6870 0.6780 1.9410 0.7020 ;
      RECT 1.3430 0.4600 1.3930 0.5020 ;
      RECT 1.0230 0.4100 1.3930 0.4600 ;
      RECT 1.0230 1.0200 1.7000 1.0700 ;
      RECT 1.6500 0.7520 1.7000 1.0200 ;
      RECT 1.6500 0.7280 1.7370 0.7520 ;
      RECT 1.6870 0.5520 1.7370 0.6780 ;
      RECT 1.3430 0.5020 1.7370 0.5520 ;
      RECT 0.8870 0.3100 1.5450 0.3600 ;
      RECT 1.4950 0.3600 1.5450 0.3920 ;
      RECT 0.8870 0.3600 0.9370 0.3920 ;
      RECT 5.6590 0.8660 5.8080 0.9160 ;
      RECT 5.7580 0.9160 5.8080 0.9670 ;
      RECT 5.7580 0.9670 5.8930 1.0170 ;
      RECT 6.8390 0.6130 7.2610 0.6630 ;
      RECT 6.8390 0.6630 6.8890 0.7590 ;
      RECT 6.3590 0.7590 6.8890 0.8090 ;
      RECT 6.3590 0.8090 6.4090 1.3010 ;
      RECT 6.3590 0.5500 6.4090 0.7590 ;
      RECT 6.1310 0.5000 6.4090 0.5500 ;
      RECT 6.1310 0.5500 6.1810 0.6790 ;
      RECT 6.6630 0.8090 6.7130 1.3010 ;
      RECT 1.9910 0.6280 2.2450 0.6520 ;
      RECT 1.9520 0.6020 2.2450 0.6280 ;
      RECT 1.9910 0.6520 2.0410 0.7780 ;
      RECT 1.9520 0.5780 2.0410 0.6020 ;
      RECT 1.9520 0.7780 2.0410 0.8280 ;
      RECT 1.9520 0.3190 2.0020 0.5780 ;
      RECT 1.9520 0.8280 2.0020 1.0760 ;
      RECT 8.4710 0.7090 9.0090 0.7590 ;
      RECT 5.2010 1.5200 8.1730 1.5700 ;
      RECT 4.6710 0.4880 5.2330 0.5380 ;
      RECT 5.1830 0.5380 5.2330 1.0200 ;
      RECT 4.6870 1.0200 5.2330 1.0700 ;
      RECT 4.4230 0.7880 4.4730 1.1200 ;
      RECT 3.3740 0.7380 4.4750 0.7880 ;
      RECT 4.2310 0.5050 4.2810 0.7380 ;
      RECT 4.6870 1.0700 4.7370 1.1200 ;
      RECT 3.9110 1.1200 4.7370 1.1700 ;
      RECT 9.0550 0.6270 9.1450 0.6770 ;
      RECT 9.0950 0.6770 9.1450 0.7680 ;
      RECT 9.0550 0.3930 9.1450 0.4430 ;
      RECT 9.0950 0.1260 9.1450 0.3930 ;
      RECT 9.0550 0.5120 9.1050 0.6270 ;
      RECT 8.8510 0.4620 9.1050 0.5120 ;
      RECT 9.0550 0.4430 9.1050 0.4620 ;
      RECT 2.9220 0.0940 3.3150 0.1440 ;
      RECT 4.4430 1.5200 5.1330 1.5700 ;
      RECT 4.8980 0.6130 5.1330 0.6630 ;
      RECT 5.4470 0.8670 5.5890 0.9170 ;
      RECT 5.4470 0.6630 5.4970 0.8670 ;
      RECT 5.4470 0.6130 5.8930 0.6630 ;
      RECT 4.5350 0.9200 4.9650 0.9700 ;
      RECT 4.9150 0.8310 4.9650 0.9200 ;
      RECT 4.5350 0.9700 4.5850 1.0340 ;
      RECT 4.5350 0.5050 4.5850 0.9200 ;
      RECT 4.2910 1.4200 5.5970 1.4700 ;
      RECT 3.3030 1.1900 3.6890 1.2400 ;
      RECT 5.8800 1.2870 6.2730 1.3370 ;
      RECT 3.2270 1.3890 3.7650 1.4390 ;
      RECT 5.1470 0.1880 5.7410 0.2380 ;
      RECT 5.1470 0.2380 5.1970 0.2880 ;
      RECT 4.5060 0.2880 5.1970 0.3380 ;
      RECT 4.1190 0.4550 4.1690 0.6130 ;
      RECT 3.6830 0.6130 4.1690 0.6630 ;
      RECT 4.5060 0.3380 4.5560 0.4050 ;
      RECT 4.1190 0.4050 4.5560 0.4550 ;
      RECT 2.6190 1.5240 3.9170 1.5740 ;
      RECT 7.1790 1.1990 8.4770 1.2490 ;
      RECT 8.4710 0.1320 8.7050 0.1820 ;
      RECT 7.7270 1.0820 8.1760 1.1320 ;
      RECT 7.7270 0.6770 7.7770 1.0820 ;
      RECT 7.6870 0.6270 7.7770 0.6770 ;
      RECT 7.6870 0.4770 7.7370 0.6270 ;
      RECT 7.6870 0.4270 7.7770 0.4770 ;
      RECT 7.7270 0.1260 7.7770 0.4270 ;
      RECT 7.7870 0.5270 8.3850 0.5770 ;
      RECT 8.0310 0.5770 8.0810 0.8780 ;
      RECT 8.0310 0.1260 8.0810 0.5270 ;
      RECT 8.3350 0.5770 8.3850 0.7700 ;
      RECT 8.3350 0.3480 8.3850 0.5270 ;
      RECT 0.7190 0.5100 1.2570 0.5600 ;
      RECT 1.1750 1.1330 1.5610 1.1830 ;
      RECT 0.7190 0.9410 0.9530 0.9910 ;
      RECT 8.6990 1.0970 9.2370 1.1470 ;
      RECT 8.1670 0.2480 9.0090 0.2980 ;
      RECT 2.8630 0.7130 2.9890 0.7630 ;
      RECT 2.8630 0.7630 2.9130 1.0330 ;
      RECT 2.9390 0.5630 2.9890 0.7130 ;
      RECT 2.8470 0.5130 2.9890 0.5630 ;
      RECT 4.8230 0.3880 5.4970 0.4380 ;
      RECT 5.4470 0.4380 5.4970 0.5630 ;
      RECT 5.4470 0.2970 5.4970 0.3880 ;
      RECT 5.2950 0.9670 5.5130 1.0170 ;
      RECT 5.2950 0.4380 5.3450 0.9670 ;
      RECT 5.2950 1.0170 5.3450 1.1200 ;
      RECT 5.2950 1.1700 5.3450 1.2700 ;
      RECT 4.8230 1.1200 5.3450 1.1700 ;
      RECT 4.2130 0.8580 4.3730 0.9080 ;
      RECT 4.2130 0.9080 4.2630 0.9680 ;
      RECT 3.6830 0.9680 4.2630 1.0180 ;
      RECT 1.4520 0.6020 1.6370 0.6520 ;
      RECT 0.2050 0.8410 1.5020 0.8910 ;
      RECT 1.4520 0.6520 1.5020 0.8410 ;
      RECT 0.2050 0.5260 0.2550 0.8410 ;
      RECT 0.2790 0.8910 0.3290 1.2140 ;
      RECT 0.2050 0.4760 0.3290 0.5260 ;
    LAYER PO ;
      RECT 5.8370 0.0660 5.8670 0.6910 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 3.1010 0.8400 3.1310 1.6060 ;
      RECT 5.8370 0.9390 5.8670 1.6060 ;
      RECT 5.5330 0.0660 5.5630 0.6370 ;
      RECT 3.1010 0.0660 3.1310 0.6370 ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 3.7090 0.0660 3.7390 0.6910 ;
      RECT 5.0770 0.0660 5.1070 0.6910 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 9.4850 0.0660 9.5150 1.6060 ;
      RECT 4.7730 0.8920 4.8030 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 5.5330 0.8390 5.5630 1.6060 ;
      RECT 9.6370 0.0660 9.6670 1.6060 ;
      RECT 10.0930 0.0660 10.1230 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 9.7890 0.0660 9.8190 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 9.9410 0.0660 9.9710 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 4.7730 0.0660 4.8030 0.6910 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 3.7090 0.9390 3.7390 1.6060 ;
      RECT 7.2050 0.0670 7.2350 1.6050 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 5.0770 0.8390 5.1070 1.6060 ;
      RECT 9.3330 0.0660 9.3630 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
    LAYER NWELL ;
      RECT 7.5600 0.4910 9.5710 1.0830 ;
      RECT -0.1150 1.5430 10.3060 1.7730 ;
      RECT -0.1150 0.6790 7.0980 1.5430 ;
      RECT 10.0310 0.6790 10.3060 1.5430 ;
  END
END RSDFFNSRASRQX1_LVT

MACRO RSDFFNSRASRQX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.336 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 10.3360 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 2.1030 1.1310 2.1530 1.6420 ;
        RECT 1.7990 1.1310 1.8490 1.6420 ;
        RECT 1.6470 1.1310 1.6970 1.6420 ;
        RECT 8.3750 1.4540 8.4250 1.6420 ;
        RECT 3.9670 1.2700 4.0170 1.6420 ;
        RECT 2.2550 1.2940 2.3050 1.6420 ;
        RECT 5.7510 1.4040 8.4250 1.4540 ;
        RECT 3.7580 1.2200 5.0570 1.2700 ;
        RECT 2.2550 1.2440 2.7770 1.2940 ;
        RECT 5.7510 1.2790 5.8010 1.4040 ;
        RECT 6.8150 0.9590 6.8650 1.4040 ;
        RECT 6.5110 0.9530 6.5610 1.4040 ;
        RECT 7.1190 1.0690 7.1690 1.4040 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 10.3360 0.0300 ;
        RECT 2.1030 0.0300 2.1530 0.3070 ;
        RECT 7.1190 0.0300 7.1690 0.2410 ;
        RECT 9.3990 0.0300 9.4490 0.4260 ;
        RECT 1.6470 0.0300 1.6970 0.4050 ;
        RECT 6.8150 0.0300 6.8650 0.2410 ;
        RECT 1.7990 0.0300 1.8490 0.4050 ;
        RECT 8.0310 0.0300 8.0810 0.4260 ;
        RECT 0.5830 0.0300 0.6330 0.5120 ;
        RECT 0.4310 0.0300 0.4810 0.4340 ;
        RECT 8.9430 0.0300 8.9930 0.1980 ;
        RECT 6.6870 0.0300 6.7370 0.2880 ;
        RECT 2.1030 0.3070 3.9770 0.3570 ;
        RECT 5.7350 0.2880 6.7370 0.3380 ;
        RECT 2.5590 0.3570 2.6090 0.5570 ;
        RECT 3.7750 0.3570 3.8250 0.5570 ;
        RECT 2.7110 0.3570 2.7610 0.5570 ;
        RECT 3.9270 0.3570 3.9770 0.5330 ;
        RECT 2.1030 0.3570 2.1530 0.4050 ;
        RECT 3.9270 0.2380 3.9770 0.3070 ;
        RECT 3.9270 0.1880 5.0570 0.2380 ;
        RECT 4.3830 0.2380 4.4330 0.3490 ;
    END
  END VSS

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.9790 0.8570 6.1350 0.9750 ;
        RECT 5.9790 0.9750 6.0290 1.0790 ;
        RECT 5.4470 1.0790 6.0290 1.1290 ;
        RECT 5.4470 1.1290 5.4970 1.3200 ;
        RECT 4.1550 1.3200 5.4970 1.3700 ;
        RECT 4.1550 1.3700 4.2050 1.4550 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4390 0.0880 6.4850 0.1380 ;
        RECT 3.4390 0.1380 3.5970 0.2100 ;
        RECT 6.4350 0.1380 6.4850 0.1700 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.9510 0.3010 7.6550 0.3510 ;
        RECT 7.5450 0.2500 7.6550 0.3010 ;
        RECT 7.5450 0.3510 7.6550 0.3600 ;
        RECT 7.6030 0.3600 7.6530 0.9690 ;
        RECT 6.9670 0.9690 7.6530 1.0190 ;
        RECT 6.9670 1.0190 7.0170 1.3270 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3770 1.4650 2.5490 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.5210 0.2490 9.6310 0.3590 ;
        RECT 9.5320 0.3590 9.5820 0.5270 ;
        RECT 9.3070 0.5270 9.5820 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6570 0.7040 4.8130 0.7310 ;
        RECT 4.6570 0.7310 5.1170 0.7810 ;
        RECT 4.7630 0.5970 4.8130 0.7040 ;
        RECT 4.6570 0.7810 4.8130 0.8150 ;
        RECT 5.0670 0.7810 5.1170 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 8.0150 0.9490 9.6330 1.0090 ;
        RECT 9.5230 0.6900 9.6330 0.9490 ;
        RECT 9.3990 0.6270 9.4490 0.9490 ;
    END
  END VDDG

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2520 1.3330 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6780 0.7250 0.7280 ;
        RECT 0.4010 0.5510 0.5110 0.6780 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 1.1610 1.0110 1.3160 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D
  OBS
    LAYER M1 ;
      RECT 0.2050 0.4760 0.3290 0.5260 ;
      RECT 0.2790 0.3160 0.3290 0.4760 ;
      RECT 3.1670 0.8540 4.0690 0.9040 ;
      RECT 3.1670 0.6130 3.2170 0.8540 ;
      RECT 3.1670 0.9040 3.2170 1.0590 ;
      RECT 3.1670 0.5630 3.3690 0.6130 ;
      RECT 3.1670 1.0590 3.5370 1.1090 ;
      RECT 3.3190 0.4070 3.3690 0.5630 ;
      RECT 3.1670 0.4130 3.2170 0.5630 ;
      RECT 3.1670 1.1090 3.2170 1.3370 ;
      RECT 5.5990 0.4000 6.6370 0.4500 ;
      RECT 6.5870 0.4500 6.6370 0.6920 ;
      RECT 5.9430 0.4500 5.9930 0.7290 ;
      RECT 5.9430 0.7290 6.3090 0.7790 ;
      RECT 6.2590 0.7790 6.3090 1.1790 ;
      RECT 5.6000 1.1790 6.3090 1.2290 ;
      RECT 5.5990 0.4500 5.6490 0.5630 ;
      RECT 5.5990 0.2970 5.6490 0.4000 ;
      RECT 5.6000 1.2290 5.6500 1.3530 ;
      RECT 6.8390 0.6130 7.4130 0.6630 ;
      RECT 6.3590 0.8090 6.4090 1.3010 ;
      RECT 6.3590 0.5500 6.4090 0.7590 ;
      RECT 6.1310 0.5000 6.4090 0.5500 ;
      RECT 6.1310 0.5500 6.1810 0.6790 ;
      RECT 6.6630 0.8090 6.7130 1.3010 ;
      RECT 6.8390 0.6630 6.8890 0.7590 ;
      RECT 6.3590 0.7590 6.8890 0.8090 ;
      RECT 5.1470 0.1880 5.7410 0.2380 ;
      RECT 5.1470 0.2380 5.1970 0.2880 ;
      RECT 4.5060 0.2880 5.1970 0.3380 ;
      RECT 4.1190 0.4550 4.1690 0.6130 ;
      RECT 3.6830 0.6130 4.1690 0.6630 ;
      RECT 4.5060 0.3380 4.5560 0.4050 ;
      RECT 4.1190 0.4050 4.5560 0.4550 ;
      RECT 3.0150 0.8130 3.1050 0.8630 ;
      RECT 3.0550 0.4620 3.1050 0.8130 ;
      RECT 3.0150 0.8630 3.0650 1.0830 ;
      RECT 2.9990 0.4120 3.1050 0.4620 ;
      RECT 2.2550 1.0830 3.0650 1.1330 ;
      RECT 3.0150 1.1330 3.0650 1.3540 ;
      RECT 2.2550 0.7520 2.3050 1.0830 ;
      RECT 2.2550 0.7020 2.3450 0.7520 ;
      RECT 2.2950 0.5510 2.3450 0.7020 ;
      RECT 2.2550 0.5010 2.3450 0.5510 ;
      RECT 2.2550 0.4070 2.3050 0.5010 ;
      RECT 2.4070 0.6130 2.8530 0.6630 ;
      RECT 2.4070 0.6630 2.4570 1.0040 ;
      RECT 2.4070 0.4130 2.4570 0.6130 ;
      RECT 8.3190 0.8200 8.8670 0.8700 ;
      RECT 1.6500 0.7020 1.9410 0.7280 ;
      RECT 1.6870 0.6780 1.9410 0.7020 ;
      RECT 1.3430 0.4600 1.3930 0.5020 ;
      RECT 1.0230 0.4100 1.3930 0.4600 ;
      RECT 1.0230 1.0200 1.7000 1.0700 ;
      RECT 1.6500 0.7520 1.7000 1.0200 ;
      RECT 1.6500 0.7280 1.7370 0.7520 ;
      RECT 1.6870 0.5520 1.7370 0.6780 ;
      RECT 1.3430 0.5020 1.7370 0.5520 ;
      RECT 0.8870 0.3100 1.5450 0.3600 ;
      RECT 1.4950 0.3600 1.5450 0.3920 ;
      RECT 0.8870 0.3600 0.9370 0.3920 ;
      RECT 5.6590 0.8660 5.8080 0.9160 ;
      RECT 5.7580 0.9160 5.8080 0.9670 ;
      RECT 5.7580 0.9670 5.8930 1.0170 ;
      RECT 1.9910 0.6280 2.2450 0.6520 ;
      RECT 1.9520 0.6020 2.2450 0.6280 ;
      RECT 1.9910 0.6520 2.0410 0.7780 ;
      RECT 1.9520 0.5780 2.0410 0.6020 ;
      RECT 1.9520 0.7780 2.0410 0.8280 ;
      RECT 1.9520 0.3190 2.0020 0.5780 ;
      RECT 1.9520 0.8280 2.0020 1.0760 ;
      RECT 8.6230 0.7090 9.1610 0.7590 ;
      RECT 8.3190 0.2480 9.1610 0.2980 ;
      RECT 5.1830 0.5380 5.2330 1.0200 ;
      RECT 4.6710 0.5110 5.2330 0.5380 ;
      RECT 4.6870 1.0200 5.2330 1.0700 ;
      RECT 4.6710 0.4880 5.2320 0.5110 ;
      RECT 4.4230 0.7880 4.4730 1.1200 ;
      RECT 3.3740 0.7380 4.4750 0.7880 ;
      RECT 4.2310 0.5050 4.2810 0.7380 ;
      RECT 4.6870 1.0700 4.7370 1.1200 ;
      RECT 3.9110 1.1200 4.7370 1.1700 ;
      RECT 5.2010 1.5200 8.3250 1.5700 ;
      RECT 9.2470 0.6770 9.2970 0.7680 ;
      RECT 9.2070 0.4270 9.2970 0.4620 ;
      RECT 9.2470 0.1260 9.2970 0.4270 ;
      RECT 9.2070 0.6270 9.2970 0.6770 ;
      RECT 9.2070 0.5120 9.2570 0.6270 ;
      RECT 9.0030 0.4770 9.2570 0.5120 ;
      RECT 9.0030 0.4620 9.2970 0.4770 ;
      RECT 2.9220 0.0940 3.3150 0.1440 ;
      RECT 4.4430 1.5200 5.1330 1.5700 ;
      RECT 4.8980 0.6130 5.1330 0.6630 ;
      RECT 5.4470 0.8670 5.5890 0.9170 ;
      RECT 5.4470 0.6630 5.4970 0.8670 ;
      RECT 5.4470 0.6130 5.8930 0.6630 ;
      RECT 4.5350 0.9200 4.9650 0.9700 ;
      RECT 4.9150 0.8310 4.9650 0.9200 ;
      RECT 4.5350 0.9700 4.5850 1.0340 ;
      RECT 4.5350 0.5050 4.5850 0.9200 ;
      RECT 4.2910 1.4200 5.5970 1.4700 ;
      RECT 3.3030 1.1900 3.6890 1.2400 ;
      RECT 5.8800 1.2870 6.2730 1.3370 ;
      RECT 3.2270 1.3890 3.7650 1.4390 ;
      RECT 2.6190 1.5240 3.9170 1.5740 ;
      RECT 7.3310 1.1990 8.6290 1.2490 ;
      RECT 7.9390 0.5270 8.5370 0.5770 ;
      RECT 8.4870 0.5770 8.5370 0.7700 ;
      RECT 8.4870 0.3480 8.5370 0.5270 ;
      RECT 8.1830 0.5770 8.2330 0.8870 ;
      RECT 8.1830 0.1260 8.2330 0.5270 ;
      RECT 8.6230 0.1320 8.8570 0.1820 ;
      RECT 7.8790 1.0770 8.3280 1.1270 ;
      RECT 7.8790 0.6770 7.9290 1.0770 ;
      RECT 7.8390 0.6270 7.9290 0.6770 ;
      RECT 7.8390 0.4770 7.8890 0.6270 ;
      RECT 7.8390 0.4270 7.9290 0.4770 ;
      RECT 7.8790 0.1260 7.9290 0.4270 ;
      RECT 0.7190 0.5100 1.2570 0.5600 ;
      RECT 1.1750 1.1330 1.5610 1.1830 ;
      RECT 0.7190 0.9410 0.9530 0.9910 ;
      RECT 8.8510 1.1050 9.3890 1.1550 ;
      RECT 2.8630 0.7130 2.9890 0.7630 ;
      RECT 2.8630 0.7630 2.9130 1.0330 ;
      RECT 2.9390 0.5630 2.9890 0.7130 ;
      RECT 2.8470 0.5130 2.9890 0.5630 ;
      RECT 4.8230 0.3880 5.4970 0.4380 ;
      RECT 5.4470 0.4380 5.4970 0.5630 ;
      RECT 5.4470 0.2970 5.4970 0.3880 ;
      RECT 5.2950 0.9670 5.5130 1.0170 ;
      RECT 5.2950 0.4380 5.3450 0.9670 ;
      RECT 5.2950 1.0170 5.3450 1.1200 ;
      RECT 5.2950 1.1700 5.3450 1.2700 ;
      RECT 4.8230 1.1200 5.3450 1.1700 ;
      RECT 4.2130 0.8580 4.3730 0.9080 ;
      RECT 4.2130 0.9080 4.2630 0.9680 ;
      RECT 3.6830 0.9680 4.2630 1.0180 ;
      RECT 1.4520 0.6020 1.6370 0.6520 ;
      RECT 0.2050 0.8410 1.5020 0.8910 ;
      RECT 1.4520 0.6520 1.5020 0.8410 ;
      RECT 0.2050 0.5260 0.2550 0.8410 ;
      RECT 0.2790 0.8910 0.3290 1.2140 ;
    LAYER PO ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 5.8370 0.0660 5.8670 0.6910 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 3.1010 0.8400 3.1310 1.6060 ;
      RECT 5.8370 0.9390 5.8670 1.6060 ;
      RECT 5.5330 0.0660 5.5630 0.6370 ;
      RECT 3.1010 0.0660 3.1310 0.6370 ;
      RECT 3.7090 0.0660 3.7390 0.6910 ;
      RECT 9.3330 0.0660 9.3630 1.6060 ;
      RECT 5.0770 0.0660 5.1070 0.6910 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 9.6370 0.0660 9.6670 1.6060 ;
      RECT 4.7730 0.8920 4.8030 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 5.5330 0.8390 5.5630 1.6060 ;
      RECT 9.7890 0.0660 9.8190 1.6060 ;
      RECT 10.2450 0.0660 10.2750 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 9.9410 0.0660 9.9710 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 10.0930 0.0660 10.1230 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 4.7730 0.0660 4.8030 0.6910 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 3.7090 0.9390 3.7390 1.6060 ;
      RECT 7.3570 0.0670 7.3870 1.6050 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 5.0770 0.8390 5.1070 1.6060 ;
      RECT 9.4850 0.0660 9.5150 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
    LAYER NWELL ;
      RECT 7.7120 0.4910 9.7230 1.0830 ;
      RECT -0.1150 1.5430 10.4580 1.7730 ;
      RECT -0.1150 0.6790 7.2500 1.5430 ;
      RECT 10.1830 0.6790 10.4580 1.5430 ;
  END
END RSDFFNSRASRQX2_LVT

MACRO RSDFFNSRASRX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.336 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 10.3360 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 2.1030 1.1310 2.1530 1.6420 ;
        RECT 1.7990 1.1310 1.8490 1.6420 ;
        RECT 1.6470 1.1310 1.6970 1.6420 ;
        RECT 8.3750 1.4540 8.4250 1.6420 ;
        RECT 3.9670 1.2700 4.0170 1.6420 ;
        RECT 2.2550 1.2940 2.3050 1.6420 ;
        RECT 5.7510 1.4040 8.4250 1.4540 ;
        RECT 3.7580 1.2200 5.0570 1.2700 ;
        RECT 2.2550 1.2440 2.7770 1.2940 ;
        RECT 5.7510 1.2790 5.8010 1.4040 ;
        RECT 6.9670 0.9590 7.0170 1.4040 ;
        RECT 6.5110 0.9530 6.5610 1.4040 ;
    END
  END VDD

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.8150 0.4010 7.5150 0.4510 ;
        RECT 6.8150 0.1570 6.8650 0.4010 ;
        RECT 7.3930 0.4510 7.5150 0.5380 ;
        RECT 7.4650 0.5380 7.5150 0.8590 ;
        RECT 6.8150 0.8590 7.5150 0.9090 ;
        RECT 6.8150 0.9090 6.8650 1.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.1190 0.9690 7.6530 1.0190 ;
        RECT 7.6030 0.3510 7.6530 0.9690 ;
        RECT 7.1190 1.0190 7.3510 1.1290 ;
        RECT 7.1030 0.3010 7.6530 0.3510 ;
        RECT 7.1190 1.1290 7.1690 1.3270 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 10.3360 0.0300 ;
        RECT 2.1030 0.0300 2.1530 0.3070 ;
        RECT 9.3990 0.0300 9.4490 0.4260 ;
        RECT 1.6470 0.0300 1.6970 0.4050 ;
        RECT 6.9670 0.0300 7.0170 0.2410 ;
        RECT 1.7990 0.0300 1.8490 0.4050 ;
        RECT 8.0310 0.0300 8.0810 0.4260 ;
        RECT 0.5830 0.0300 0.6330 0.5120 ;
        RECT 0.4310 0.0300 0.4810 0.4340 ;
        RECT 8.9430 0.0300 8.9930 0.1980 ;
        RECT 6.6870 0.0300 6.7370 0.2930 ;
        RECT 2.1030 0.3070 3.9770 0.3570 ;
        RECT 5.7350 0.2930 6.7370 0.3400 ;
        RECT 2.5590 0.3570 2.6090 0.5570 ;
        RECT 3.7750 0.3570 3.8250 0.5570 ;
        RECT 2.7110 0.3570 2.7610 0.5570 ;
        RECT 3.9270 0.3570 3.9770 0.5330 ;
        RECT 2.1030 0.3570 2.1530 0.4050 ;
        RECT 3.9270 0.2440 3.9770 0.3070 ;
        RECT 5.7350 0.3400 6.7120 0.3430 ;
        RECT 3.9270 0.1940 5.0570 0.2440 ;
        RECT 4.3830 0.2440 4.4330 0.3490 ;
    END
  END VSS

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.9790 0.8570 6.1350 0.9750 ;
        RECT 5.9790 0.9750 6.0290 1.0790 ;
        RECT 5.4470 1.0790 6.0290 1.1290 ;
        RECT 5.4470 1.1290 5.4970 1.3200 ;
        RECT 4.1550 1.3200 5.4970 1.3700 ;
        RECT 4.1550 1.3700 4.2050 1.4550 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4390 0.0880 6.5210 0.1380 ;
        RECT 3.4390 0.1380 3.5970 0.2100 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3770 1.4650 2.5490 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.5210 0.2490 9.6310 0.3590 ;
        RECT 9.5320 0.3590 9.5820 0.5270 ;
        RECT 9.3070 0.5270 9.5820 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6570 0.7050 4.8130 0.7310 ;
        RECT 4.6570 0.7310 5.1170 0.7810 ;
        RECT 4.7630 0.5970 4.8130 0.7050 ;
        RECT 4.6570 0.7810 4.8130 0.8150 ;
        RECT 5.0670 0.7810 5.1170 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 8.0150 0.9500 9.6330 1.0100 ;
        RECT 9.5230 0.6900 9.6330 0.9500 ;
        RECT 9.3990 0.6270 9.4490 0.9500 ;
    END
  END VDDG

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2520 1.3330 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6780 0.7250 0.7280 ;
        RECT 0.4010 0.5510 0.5110 0.6780 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 1.1610 1.0110 1.3160 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D
  OBS
    LAYER M1 ;
      RECT 5.2950 1.0170 5.3450 1.1200 ;
      RECT 5.2950 1.1700 5.3450 1.2700 ;
      RECT 4.8230 1.1200 5.3450 1.1700 ;
      RECT 4.2130 0.8580 4.3730 0.9080 ;
      RECT 4.2130 0.9080 4.2630 0.9680 ;
      RECT 3.6830 0.9680 4.2630 1.0180 ;
      RECT 1.4520 0.6020 1.6370 0.6520 ;
      RECT 0.2050 0.8410 1.5020 0.8910 ;
      RECT 1.4520 0.6520 1.5020 0.8410 ;
      RECT 0.2050 0.5260 0.2550 0.8410 ;
      RECT 0.2790 0.8910 0.3290 1.2140 ;
      RECT 0.2050 0.4760 0.3290 0.5260 ;
      RECT 0.2790 0.3160 0.3290 0.4760 ;
      RECT 3.1670 0.8540 4.0690 0.9040 ;
      RECT 3.1670 0.6130 3.2170 0.8540 ;
      RECT 3.1670 0.9040 3.2170 1.0590 ;
      RECT 3.1670 0.5630 3.3690 0.6130 ;
      RECT 3.1670 1.0590 3.5370 1.1090 ;
      RECT 3.3190 0.4070 3.3690 0.5630 ;
      RECT 3.1670 0.4130 3.2170 0.5630 ;
      RECT 3.1670 1.1090 3.2170 1.3370 ;
      RECT 6.5870 0.6320 6.9410 0.6820 ;
      RECT 6.8910 0.5970 6.9410 0.6320 ;
      RECT 6.2590 0.7790 6.3090 1.1790 ;
      RECT 5.9430 0.7290 6.3090 0.7790 ;
      RECT 5.9430 0.4500 5.9930 0.7290 ;
      RECT 5.5990 0.4000 6.6370 0.4500 ;
      RECT 6.5870 0.4500 6.6370 0.6320 ;
      RECT 5.6000 1.1790 6.3090 1.2290 ;
      RECT 5.6000 1.2290 5.6500 1.3530 ;
      RECT 5.5990 0.4500 5.6490 0.5630 ;
      RECT 5.5990 0.2970 5.6490 0.4000 ;
      RECT 5.1470 0.1880 5.7410 0.2380 ;
      RECT 5.1470 0.2380 5.1970 0.2940 ;
      RECT 4.5060 0.2940 5.1970 0.3440 ;
      RECT 4.1190 0.4550 4.1690 0.6130 ;
      RECT 3.6830 0.6130 4.1690 0.6630 ;
      RECT 4.5060 0.3440 4.5560 0.4050 ;
      RECT 4.1190 0.4050 4.5560 0.4550 ;
      RECT 6.9910 0.6130 7.4130 0.6630 ;
      RECT 6.3590 0.8090 6.4090 1.3010 ;
      RECT 6.3590 0.5500 6.4090 0.7590 ;
      RECT 6.1310 0.5000 6.4090 0.5500 ;
      RECT 6.1310 0.5500 6.1810 0.6790 ;
      RECT 6.6630 0.8090 6.7130 1.3010 ;
      RECT 6.9910 0.6630 7.0410 0.7590 ;
      RECT 6.3590 0.7590 7.0410 0.8090 ;
      RECT 3.0150 0.8130 3.1050 0.8630 ;
      RECT 3.0550 0.4620 3.1050 0.8130 ;
      RECT 3.0150 0.8630 3.0650 1.0830 ;
      RECT 2.9990 0.4120 3.1050 0.4620 ;
      RECT 2.2550 1.0830 3.0650 1.1330 ;
      RECT 3.0150 1.1330 3.0650 1.3540 ;
      RECT 2.2550 0.7520 2.3050 1.0830 ;
      RECT 2.2550 0.7020 2.3450 0.7520 ;
      RECT 2.2950 0.5510 2.3450 0.7020 ;
      RECT 2.2550 0.5010 2.3450 0.5510 ;
      RECT 2.2550 0.4070 2.3050 0.5010 ;
      RECT 2.4070 0.6130 2.8530 0.6630 ;
      RECT 2.4070 0.6630 2.4570 1.0040 ;
      RECT 2.4070 0.4130 2.4570 0.6130 ;
      RECT 8.3190 0.8200 8.8670 0.8700 ;
      RECT 1.6500 0.7020 1.9410 0.7280 ;
      RECT 1.6870 0.6780 1.9410 0.7020 ;
      RECT 1.3430 0.4600 1.3930 0.5020 ;
      RECT 1.0230 0.4100 1.3930 0.4600 ;
      RECT 1.0230 1.0200 1.7000 1.0700 ;
      RECT 1.6500 0.7520 1.7000 1.0200 ;
      RECT 1.6500 0.7280 1.7370 0.7520 ;
      RECT 1.6870 0.5520 1.7370 0.6780 ;
      RECT 1.3430 0.5020 1.7370 0.5520 ;
      RECT 0.8870 0.3100 1.5450 0.3600 ;
      RECT 1.4950 0.3600 1.5450 0.3920 ;
      RECT 0.8870 0.3600 0.9370 0.3920 ;
      RECT 5.6590 0.8660 5.8080 0.9160 ;
      RECT 5.7580 0.9160 5.8080 0.9670 ;
      RECT 5.7580 0.9670 5.8930 1.0170 ;
      RECT 1.9910 0.6280 2.2450 0.6520 ;
      RECT 1.9520 0.6020 2.2450 0.6280 ;
      RECT 1.9910 0.6520 2.0410 0.7780 ;
      RECT 1.9520 0.5780 2.0410 0.6020 ;
      RECT 1.9520 0.7780 2.0410 0.8280 ;
      RECT 1.9520 0.3190 2.0020 0.5780 ;
      RECT 1.9520 0.8280 2.0020 1.0760 ;
      RECT 8.6230 0.7090 9.1610 0.7590 ;
      RECT 4.6710 0.4940 5.2320 0.5170 ;
      RECT 4.6710 0.5170 5.2330 0.5440 ;
      RECT 5.1830 0.5440 5.2330 1.0200 ;
      RECT 4.6870 1.0200 5.2330 1.0700 ;
      RECT 4.4230 0.7880 4.4730 1.1200 ;
      RECT 3.3740 0.7380 4.4750 0.7880 ;
      RECT 4.2310 0.5050 4.2810 0.7380 ;
      RECT 4.6870 1.0700 4.7370 1.1200 ;
      RECT 3.9110 1.1200 4.7370 1.1700 ;
      RECT 5.2010 1.5200 8.3250 1.5700 ;
      RECT 9.2470 0.6770 9.2970 0.7680 ;
      RECT 9.2070 0.4270 9.2970 0.4620 ;
      RECT 9.2470 0.1260 9.2970 0.4270 ;
      RECT 9.2070 0.6270 9.2970 0.6770 ;
      RECT 9.2070 0.5120 9.2570 0.6270 ;
      RECT 9.0030 0.4770 9.2570 0.5120 ;
      RECT 9.0030 0.4620 9.2970 0.4770 ;
      RECT 2.9220 0.0940 3.3150 0.1440 ;
      RECT 4.4430 1.5200 5.1330 1.5700 ;
      RECT 4.8980 0.6130 5.1330 0.6630 ;
      RECT 5.4470 0.8670 5.5890 0.9170 ;
      RECT 5.4470 0.6630 5.4970 0.8670 ;
      RECT 5.4470 0.6130 5.8930 0.6630 ;
      RECT 4.5350 0.9200 4.9650 0.9700 ;
      RECT 4.9150 0.8310 4.9650 0.9200 ;
      RECT 4.5350 0.9700 4.5850 1.0340 ;
      RECT 4.5350 0.5050 4.5850 0.9200 ;
      RECT 4.2910 1.4200 5.5970 1.4700 ;
      RECT 3.3030 1.1900 3.6890 1.2400 ;
      RECT 5.8800 1.2870 6.2730 1.3370 ;
      RECT 3.2270 1.3890 3.7650 1.4390 ;
      RECT 2.6190 1.5240 3.9170 1.5740 ;
      RECT 7.3310 1.2140 8.6290 1.2640 ;
      RECT 7.9390 0.5270 8.5370 0.5770 ;
      RECT 8.4870 0.5770 8.5370 0.7700 ;
      RECT 8.4870 0.3480 8.5370 0.5270 ;
      RECT 8.1830 0.5770 8.2330 0.8870 ;
      RECT 8.1830 0.1260 8.2330 0.5270 ;
      RECT 8.6230 0.1320 8.8570 0.1820 ;
      RECT 7.8790 1.1070 8.3280 1.1570 ;
      RECT 7.8790 0.6770 7.9290 1.1070 ;
      RECT 7.8390 0.6270 7.9290 0.6770 ;
      RECT 7.8390 0.4770 7.8890 0.6270 ;
      RECT 7.8390 0.4270 7.9290 0.4770 ;
      RECT 7.8790 0.1260 7.9290 0.4270 ;
      RECT 0.7190 0.5100 1.2570 0.5600 ;
      RECT 1.1750 1.1330 1.5610 1.1830 ;
      RECT 0.7190 0.9410 0.9530 0.9910 ;
      RECT 8.8510 1.1270 9.3890 1.1770 ;
      RECT 8.3190 0.2480 9.1610 0.2980 ;
      RECT 2.8630 0.7130 2.9890 0.7630 ;
      RECT 2.8630 0.7630 2.9130 1.0330 ;
      RECT 2.9390 0.5630 2.9890 0.7130 ;
      RECT 2.8470 0.5130 2.9890 0.5630 ;
      RECT 4.8230 0.3940 5.4970 0.4440 ;
      RECT 5.4470 0.4440 5.4970 0.5630 ;
      RECT 5.4470 0.2970 5.4970 0.3940 ;
      RECT 5.2950 0.9670 5.5130 1.0170 ;
      RECT 5.2950 0.4440 5.3450 0.9670 ;
    LAYER PO ;
      RECT 5.0770 0.8390 5.1070 1.6060 ;
      RECT 9.4850 0.0660 9.5150 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 5.8370 0.0660 5.8670 0.6910 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 3.1010 0.8400 3.1310 1.6060 ;
      RECT 5.8370 0.9390 5.8670 1.6060 ;
      RECT 5.5330 0.0660 5.5630 0.6370 ;
      RECT 3.1010 0.0660 3.1310 0.6370 ;
      RECT 9.3330 0.0660 9.3630 1.6060 ;
      RECT 3.7090 0.0660 3.7390 0.6910 ;
      RECT 5.0770 0.0660 5.1070 0.6910 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 9.6370 0.0660 9.6670 1.6060 ;
      RECT 4.7730 0.8920 4.8030 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 5.5330 0.8390 5.5630 1.6060 ;
      RECT 9.7890 0.0660 9.8190 1.6060 ;
      RECT 10.2450 0.0660 10.2750 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 9.9410 0.0660 9.9710 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 10.0930 0.0660 10.1230 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 4.7730 0.0660 4.8030 0.6910 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 3.7090 0.9390 3.7390 1.6060 ;
      RECT 7.3570 0.0670 7.3870 1.6050 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
    LAYER NWELL ;
      RECT 7.7120 0.4910 9.7230 1.0830 ;
      RECT -0.1150 1.5430 10.4580 1.7730 ;
      RECT -0.1150 0.6790 7.2500 1.5430 ;
      RECT 10.1830 0.6790 10.4580 1.5430 ;
  END
END RSDFFNSRASRX1_LVT

MACRO RSDFFNSRASRX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.64 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 10.6400 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 1.6470 1.1310 1.6970 1.6420 ;
        RECT 2.1030 1.1310 2.1530 1.6420 ;
        RECT 1.7990 1.1310 1.8490 1.6420 ;
        RECT 2.2550 1.2940 2.3050 1.6420 ;
        RECT 3.9670 1.2700 4.0170 1.6420 ;
        RECT 8.6790 1.4540 8.7290 1.6420 ;
        RECT 2.2550 1.2440 2.7770 1.2940 ;
        RECT 3.7580 1.2200 5.0570 1.2700 ;
        RECT 5.7510 1.4040 8.7290 1.4540 ;
        RECT 5.7510 1.2790 5.8010 1.4040 ;
        RECT 7.1190 0.9610 7.1690 1.4040 ;
        RECT 6.5110 0.9530 6.5610 1.4040 ;
        RECT 7.4230 1.0530 7.4730 1.4040 ;
        RECT 6.8150 0.9130 6.8650 1.4040 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 10.6400 0.0300 ;
        RECT 2.1030 0.0300 2.1530 0.3070 ;
        RECT 1.6470 0.0300 1.6970 0.4050 ;
        RECT 0.5830 0.0300 0.6330 0.5120 ;
        RECT 0.4310 0.0300 0.4810 0.4340 ;
        RECT 1.7990 0.0300 1.8490 0.4050 ;
        RECT 6.8150 0.0300 6.8650 0.4090 ;
        RECT 7.1190 0.0300 7.1690 0.3200 ;
        RECT 8.3350 0.0300 8.3850 0.4260 ;
        RECT 7.4230 0.0300 7.4730 0.2210 ;
        RECT 9.7030 0.0300 9.7530 0.4260 ;
        RECT 9.2470 0.0300 9.2970 0.1980 ;
        RECT 6.6870 0.0300 6.7370 0.2880 ;
        RECT 2.1030 0.3070 3.9770 0.3570 ;
        RECT 5.7350 0.2880 6.7370 0.3380 ;
        RECT 3.7750 0.3570 3.8250 0.5570 ;
        RECT 2.5590 0.3570 2.6090 0.5570 ;
        RECT 2.7110 0.3570 2.7610 0.5570 ;
        RECT 3.9270 0.3570 3.9770 0.5330 ;
        RECT 2.1030 0.3570 2.1530 0.4050 ;
        RECT 3.9270 0.2380 3.9770 0.3070 ;
        RECT 3.9270 0.1880 5.0570 0.2380 ;
        RECT 4.3830 0.2380 4.4330 0.3490 ;
    END
  END VSS

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.9790 0.8570 6.1350 0.9750 ;
        RECT 5.9790 0.9750 6.0290 1.0790 ;
        RECT 5.4470 1.0790 6.0290 1.1290 ;
        RECT 5.4470 1.1290 5.4970 1.3200 ;
        RECT 4.1550 1.3200 5.4970 1.3700 ;
        RECT 4.1550 1.3700 4.2050 1.4550 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.5470 0.0880 6.4850 0.0970 ;
        RECT 3.4390 0.0970 6.4850 0.1380 ;
        RECT 3.4390 0.1380 3.5970 0.2100 ;
        RECT 6.4350 0.1380 6.4850 0.1700 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.9670 0.1490 7.0170 0.4020 ;
        RECT 6.9670 0.4020 7.8190 0.4520 ;
        RECT 7.6970 0.4520 7.8190 0.5120 ;
        RECT 7.7690 0.5120 7.8190 0.8420 ;
        RECT 6.9670 0.8420 7.8190 0.8920 ;
        RECT 6.9670 0.8920 7.0170 1.3190 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3770 1.4650 2.5490 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.8250 0.2490 9.9350 0.3590 ;
        RECT 9.8360 0.3590 9.8860 0.5270 ;
        RECT 9.6110 0.5270 9.8860 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.7630 0.5970 4.8130 0.7050 ;
        RECT 4.6570 0.7050 4.8130 0.7310 ;
        RECT 4.6570 0.7310 5.1170 0.7810 ;
        RECT 4.6570 0.7810 4.8130 0.8150 ;
        RECT 5.0670 0.7810 5.1170 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.2710 0.1490 7.3210 0.2710 ;
        RECT 7.2710 0.2710 7.9690 0.3210 ;
        RECT 7.8480 0.3210 7.9690 0.3600 ;
        RECT 7.8480 0.2500 7.9690 0.2710 ;
        RECT 7.9190 0.3600 7.9690 0.9420 ;
        RECT 7.8480 0.2480 7.9610 0.2500 ;
        RECT 7.2710 0.9420 7.9690 0.9920 ;
        RECT 7.2710 0.9920 7.3210 1.3270 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 8.3190 0.9490 9.9370 1.0090 ;
        RECT 9.8270 0.6900 9.9370 0.9490 ;
        RECT 9.7030 0.6270 9.7530 0.9490 ;
    END
  END VDDG

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2520 1.3330 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6780 0.7250 0.7280 ;
        RECT 0.4010 0.5510 0.5110 0.6780 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 1.1610 1.0110 1.3160 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D
  OBS
    LAYER M1 ;
      RECT 0.2050 0.8410 1.5020 0.8910 ;
      RECT 1.4520 0.6520 1.5020 0.8410 ;
      RECT 0.2050 0.5260 0.2550 0.8410 ;
      RECT 0.2790 0.8910 0.3290 1.2140 ;
      RECT 0.2050 0.4760 0.3290 0.5260 ;
      RECT 0.2790 0.3160 0.3290 0.4760 ;
      RECT 0.8870 0.3100 1.5450 0.3600 ;
      RECT 1.4950 0.3600 1.5450 0.3920 ;
      RECT 0.8870 0.3600 0.9370 0.3920 ;
      RECT 1.6870 0.6780 1.9410 0.7020 ;
      RECT 1.6500 0.7020 1.9410 0.7280 ;
      RECT 1.3430 0.4600 1.3930 0.5020 ;
      RECT 1.0230 0.4100 1.3930 0.4600 ;
      RECT 1.3430 0.5020 1.7370 0.5520 ;
      RECT 1.6870 0.5520 1.7370 0.6780 ;
      RECT 1.6500 0.7280 1.7370 0.7520 ;
      RECT 1.6500 0.7520 1.7000 1.0200 ;
      RECT 1.0230 1.0200 1.7000 1.0700 ;
      RECT 0.7190 0.5100 1.2570 0.5600 ;
      RECT 3.1670 0.8540 4.0690 0.9040 ;
      RECT 3.1670 0.9040 3.2170 1.0590 ;
      RECT 3.1670 1.0590 3.5370 1.1090 ;
      RECT 3.1670 0.6130 3.2170 0.8540 ;
      RECT 3.1670 1.1090 3.2170 1.3370 ;
      RECT 3.1670 0.5630 3.3690 0.6130 ;
      RECT 3.3190 0.4070 3.3690 0.5630 ;
      RECT 3.1670 0.4130 3.2170 0.5630 ;
      RECT 1.9910 0.6280 2.2450 0.6520 ;
      RECT 1.9520 0.6020 2.2450 0.6280 ;
      RECT 1.9910 0.6520 2.0410 0.7780 ;
      RECT 1.9520 0.5780 2.0410 0.6020 ;
      RECT 1.9520 0.7780 2.0410 0.8280 ;
      RECT 1.9520 0.3190 2.0020 0.5780 ;
      RECT 1.9520 0.8280 2.0020 1.0760 ;
      RECT 2.8470 0.5130 2.9890 0.5630 ;
      RECT 2.9390 0.5630 2.9890 0.7130 ;
      RECT 2.8630 0.7130 2.9890 0.7630 ;
      RECT 2.8630 0.7630 2.9130 1.0330 ;
      RECT 2.9990 0.4120 3.1050 0.4620 ;
      RECT 3.0550 0.4620 3.1050 0.8130 ;
      RECT 3.0150 0.8130 3.1050 0.8630 ;
      RECT 3.0150 0.8630 3.0650 1.0830 ;
      RECT 2.2550 1.0830 3.0650 1.1330 ;
      RECT 3.0150 1.1330 3.0650 1.3540 ;
      RECT 2.2550 0.7520 2.3050 1.0830 ;
      RECT 2.2550 0.7020 2.3450 0.7520 ;
      RECT 2.2950 0.5510 2.3450 0.7020 ;
      RECT 2.2550 0.5010 2.3450 0.5510 ;
      RECT 2.2550 0.4070 2.3050 0.5010 ;
      RECT 2.4070 0.6130 2.8530 0.6630 ;
      RECT 2.4070 0.6630 2.4570 1.0040 ;
      RECT 2.4070 0.4130 2.4570 0.6130 ;
      RECT 2.9220 0.0940 3.3150 0.1440 ;
      RECT 5.1470 0.1880 5.7410 0.2380 ;
      RECT 5.1470 0.2380 5.1970 0.2880 ;
      RECT 4.5060 0.2880 5.1970 0.3380 ;
      RECT 4.1190 0.4550 4.1690 0.6130 ;
      RECT 3.6830 0.6130 4.1690 0.6630 ;
      RECT 4.5060 0.3380 4.5560 0.4050 ;
      RECT 4.1190 0.4050 4.5560 0.4550 ;
      RECT 4.8230 0.3880 5.4970 0.4380 ;
      RECT 5.4470 0.4380 5.4970 0.5630 ;
      RECT 5.4470 0.2970 5.4970 0.3880 ;
      RECT 5.2950 0.9670 5.5130 1.0170 ;
      RECT 5.2950 0.4380 5.3450 0.9670 ;
      RECT 5.2950 1.0170 5.3450 1.1200 ;
      RECT 5.2950 1.1700 5.3450 1.2700 ;
      RECT 4.8230 1.1200 5.3450 1.1700 ;
      RECT 6.5870 0.6420 7.1090 0.6920 ;
      RECT 5.9430 0.4500 5.9930 0.7290 ;
      RECT 5.9430 0.7290 6.3090 0.7790 ;
      RECT 6.2590 0.7790 6.3090 1.1790 ;
      RECT 6.5870 0.4500 6.6370 0.6420 ;
      RECT 5.5990 0.4000 6.6370 0.4500 ;
      RECT 5.6000 1.1790 6.3090 1.2290 ;
      RECT 5.5990 0.4500 5.6490 0.5630 ;
      RECT 5.5990 0.2970 5.6490 0.4000 ;
      RECT 5.6000 1.2290 5.6500 1.3530 ;
      RECT 4.6710 0.4880 5.2330 0.5380 ;
      RECT 5.1830 0.5380 5.2330 1.0200 ;
      RECT 4.6870 1.0200 5.2330 1.0700 ;
      RECT 4.4230 0.7880 4.4730 1.1200 ;
      RECT 3.3740 0.7380 4.4750 0.7880 ;
      RECT 4.2310 0.5050 4.2810 0.7380 ;
      RECT 4.6870 1.0700 4.7370 1.1200 ;
      RECT 3.9110 1.1200 4.7370 1.1700 ;
      RECT 4.8980 0.6130 5.1330 0.6630 ;
      RECT 5.4470 0.6130 5.8930 0.6630 ;
      RECT 5.4470 0.6630 5.4970 0.8670 ;
      RECT 5.4470 0.8670 5.5890 0.9170 ;
      RECT 4.5350 0.9200 4.9650 0.9700 ;
      RECT 4.9150 0.8310 4.9650 0.9200 ;
      RECT 4.5350 0.9700 4.5850 1.0340 ;
      RECT 4.5350 0.5050 4.5850 0.9200 ;
      RECT 7.1590 0.6130 7.7170 0.6630 ;
      RECT 6.3590 0.7920 6.4090 1.3010 ;
      RECT 6.3590 0.5500 6.4090 0.7420 ;
      RECT 6.1310 0.5000 6.4090 0.5500 ;
      RECT 6.1310 0.5500 6.1810 0.6790 ;
      RECT 6.6630 0.7920 6.7130 1.3010 ;
      RECT 7.1590 0.6630 7.2090 0.7420 ;
      RECT 6.3590 0.7420 7.2090 0.7920 ;
      RECT 8.1830 1.0820 8.6320 1.1320 ;
      RECT 8.1830 0.6770 8.2330 1.0820 ;
      RECT 8.1430 0.6270 8.2330 0.6770 ;
      RECT 8.1430 0.4770 8.1930 0.6270 ;
      RECT 8.1430 0.4270 8.2330 0.4770 ;
      RECT 8.1830 0.1260 8.2330 0.4270 ;
      RECT 8.2430 0.5270 8.8410 0.5770 ;
      RECT 8.7910 0.5770 8.8410 0.7700 ;
      RECT 8.7910 0.3480 8.8410 0.5270 ;
      RECT 8.4870 0.5770 8.5370 0.8870 ;
      RECT 8.4870 0.1260 8.5370 0.5270 ;
      RECT 8.6230 0.2480 9.4650 0.2980 ;
      RECT 9.5510 0.6770 9.6010 0.7680 ;
      RECT 9.5110 0.4270 9.6010 0.4620 ;
      RECT 9.5510 0.1260 9.6010 0.4270 ;
      RECT 9.5110 0.6270 9.6010 0.6770 ;
      RECT 9.5110 0.5120 9.5610 0.6270 ;
      RECT 9.3070 0.4770 9.5610 0.5120 ;
      RECT 9.3070 0.4620 9.6010 0.4770 ;
      RECT 8.9270 0.1320 9.1610 0.1820 ;
      RECT 1.1750 1.1330 1.5610 1.1830 ;
      RECT 0.7190 0.9410 0.9530 0.9910 ;
      RECT 3.3030 1.1900 3.6890 1.2400 ;
      RECT 3.2270 1.3890 3.7650 1.4390 ;
      RECT 2.6190 1.5240 3.9170 1.5740 ;
      RECT 3.6830 0.9680 4.2630 1.0180 ;
      RECT 4.2130 0.9080 4.2630 0.9680 ;
      RECT 4.2130 0.8580 4.3730 0.9080 ;
      RECT 5.7580 0.9670 5.8930 1.0170 ;
      RECT 5.7580 0.9160 5.8080 0.9670 ;
      RECT 5.6590 0.8660 5.8080 0.9160 ;
      RECT 4.4430 1.5200 5.1330 1.5700 ;
      RECT 4.2910 1.4200 5.5970 1.4700 ;
      RECT 5.8800 1.2870 6.2730 1.3370 ;
      RECT 7.6350 1.2420 8.9330 1.2920 ;
      RECT 8.6230 0.8200 9.1710 0.8700 ;
      RECT 8.9270 0.7090 9.4650 0.7590 ;
      RECT 9.1550 1.1100 9.6930 1.1600 ;
      RECT 5.2010 1.5200 8.6290 1.5700 ;
      RECT 1.4520 0.6020 1.6370 0.6520 ;
    LAYER PO ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 3.7090 0.9390 3.7390 1.6060 ;
      RECT 7.6610 0.0670 7.6910 1.6050 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 9.3330 0.0660 9.3630 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 5.0770 0.8390 5.1070 1.6060 ;
      RECT 9.7890 0.0660 9.8190 1.6060 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 9.4850 0.0660 9.5150 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 5.8370 0.0660 5.8670 0.6910 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 3.1010 0.8400 3.1310 1.6060 ;
      RECT 5.8370 0.9390 5.8670 1.6060 ;
      RECT 5.5330 0.0660 5.5630 0.6370 ;
      RECT 3.7090 0.0660 3.7390 0.6910 ;
      RECT 3.1010 0.0660 3.1310 0.6370 ;
      RECT 9.6370 0.0660 9.6670 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 5.0770 0.0660 5.1070 0.6910 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 9.9410 0.0660 9.9710 1.6060 ;
      RECT 4.7730 0.8920 4.8030 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 5.5330 0.8390 5.5630 1.6060 ;
      RECT 10.0930 0.0660 10.1230 1.6060 ;
      RECT 10.5490 0.0660 10.5790 1.6060 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 10.2450 0.0660 10.2750 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 10.3970 0.0660 10.4270 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 4.7730 0.0660 4.8030 0.6910 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
    LAYER NWELL ;
      RECT 8.0160 0.4910 10.0270 1.0830 ;
      RECT -0.1150 1.5430 10.7620 1.7730 ;
      RECT -0.1150 0.6790 7.5540 1.5430 ;
      RECT 10.4870 0.6790 10.7620 1.5430 ;
  END
END RSDFFNSRASRX2_LVT

MACRO RSDFFNSRASX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.336 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3770 1.4650 2.5490 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 10.3360 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 2.1030 1.1310 2.1530 1.6420 ;
        RECT 1.7990 1.1310 1.8490 1.6420 ;
        RECT 1.6470 1.1310 1.6970 1.6420 ;
        RECT 8.3750 1.4540 8.4250 1.6420 ;
        RECT 2.2550 1.2940 2.3050 1.6420 ;
        RECT 3.9670 1.2700 4.0170 1.6420 ;
        RECT 5.7510 1.4040 8.4250 1.4540 ;
        RECT 2.2550 1.2440 2.7770 1.2940 ;
        RECT 3.7580 1.2200 5.0570 1.2700 ;
        RECT 5.7510 1.2790 5.8010 1.4040 ;
        RECT 6.9670 0.9590 7.0170 1.4040 ;
        RECT 6.5110 0.9530 6.5610 1.4040 ;
    END
  END VDD

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.8150 0.4010 7.5150 0.4510 ;
        RECT 6.8150 0.1570 6.8650 0.4010 ;
        RECT 7.3930 0.4510 7.5150 0.5380 ;
        RECT 7.4650 0.5380 7.5150 0.8590 ;
        RECT 6.8150 0.8590 7.5150 0.9090 ;
        RECT 6.8150 0.9090 6.8650 1.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.1190 0.9690 7.6530 1.0190 ;
        RECT 7.6030 0.3510 7.6530 0.9690 ;
        RECT 7.1190 1.0190 7.3510 1.1290 ;
        RECT 7.1030 0.3010 7.6530 0.3510 ;
        RECT 7.1190 1.1290 7.1690 1.3270 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 10.3360 0.0300 ;
        RECT 2.1030 0.0300 2.1530 0.3070 ;
        RECT 9.3990 0.0300 9.4490 0.4260 ;
        RECT 1.6470 0.0300 1.6970 0.4050 ;
        RECT 6.9670 0.0300 7.0170 0.2410 ;
        RECT 1.7990 0.0300 1.8490 0.4050 ;
        RECT 8.0310 0.0300 8.0810 0.4260 ;
        RECT 0.5830 0.0300 0.6330 0.5120 ;
        RECT 0.4310 0.0300 0.4810 0.4340 ;
        RECT 8.9430 0.0300 8.9930 0.1980 ;
        RECT 6.6870 0.0300 6.7370 0.2880 ;
        RECT 2.1030 0.3070 3.9770 0.3570 ;
        RECT 5.7350 0.2880 6.7370 0.3380 ;
        RECT 2.5590 0.3570 2.6090 0.5570 ;
        RECT 3.7750 0.3570 3.8250 0.5570 ;
        RECT 2.7110 0.3570 2.7610 0.5570 ;
        RECT 3.9270 0.3570 3.9770 0.5330 ;
        RECT 2.1030 0.3570 2.1530 0.4050 ;
        RECT 3.9270 0.2380 3.9770 0.3070 ;
        RECT 3.9270 0.1880 5.0570 0.2380 ;
        RECT 4.3830 0.2380 4.4330 0.3490 ;
    END
  END VSS

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.9790 0.8570 6.1350 0.9750 ;
        RECT 5.9790 0.9750 6.0290 1.0790 ;
        RECT 5.4470 1.0790 6.0290 1.1290 ;
        RECT 5.4470 1.1290 5.4970 1.3200 ;
        RECT 4.1550 1.3200 5.4970 1.3700 ;
        RECT 4.1550 1.3700 4.2050 1.4550 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.5210 0.2490 9.6310 0.3590 ;
        RECT 9.5320 0.3590 9.5820 0.5270 ;
        RECT 9.3070 0.5270 9.5820 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6570 0.7050 4.8130 0.7310 ;
        RECT 4.6570 0.7310 5.1170 0.7810 ;
        RECT 4.7630 0.5970 4.8130 0.7050 ;
        RECT 4.6570 0.7810 4.8130 0.8150 ;
        RECT 5.0670 0.7810 5.1170 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 8.0150 0.9430 9.6330 1.0030 ;
        RECT 9.5230 0.6900 9.6330 0.9430 ;
        RECT 9.3990 0.6270 9.4490 0.9430 ;
    END
  END VDDG

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2520 1.3330 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6780 0.7250 0.7280 ;
        RECT 0.4010 0.5510 0.5110 0.6780 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 1.1610 1.0110 1.3160 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D
  OBS
    LAYER M1 ;
      RECT 5.2950 0.9670 5.5130 1.0170 ;
      RECT 5.2950 0.4380 5.3450 0.9670 ;
      RECT 5.2950 1.0170 5.3450 1.1200 ;
      RECT 5.2950 1.1700 5.3450 1.2700 ;
      RECT 4.8230 1.1200 5.3450 1.1700 ;
      RECT 4.2130 0.8580 4.3730 0.9080 ;
      RECT 4.2130 0.9080 4.2630 0.9680 ;
      RECT 3.6830 0.9680 4.2630 1.0180 ;
      RECT 1.4520 0.6020 1.6370 0.6520 ;
      RECT 0.2050 0.8410 1.5020 0.8910 ;
      RECT 1.4520 0.6520 1.5020 0.8410 ;
      RECT 0.2050 0.5260 0.2550 0.8410 ;
      RECT 0.2790 0.8910 0.3290 1.2140 ;
      RECT 0.2050 0.4760 0.3290 0.5260 ;
      RECT 0.2790 0.3160 0.3290 0.4760 ;
      RECT 3.1670 0.8540 4.0690 0.9040 ;
      RECT 3.1670 0.6130 3.2170 0.8540 ;
      RECT 3.1670 0.9040 3.2170 1.0590 ;
      RECT 3.1670 0.5630 3.3690 0.6130 ;
      RECT 3.1670 1.0590 3.5370 1.1090 ;
      RECT 3.3190 0.4070 3.3690 0.5630 ;
      RECT 3.1670 0.4130 3.2170 0.5630 ;
      RECT 3.1670 1.1090 3.2170 1.3370 ;
      RECT 6.5440 0.6320 6.9410 0.6820 ;
      RECT 6.8910 0.5970 6.9410 0.6320 ;
      RECT 5.9430 0.4500 5.9930 0.7290 ;
      RECT 5.9430 0.7290 6.3090 0.7790 ;
      RECT 6.2590 0.7790 6.3090 1.1790 ;
      RECT 5.5990 0.4000 6.6370 0.4500 ;
      RECT 6.5870 0.4500 6.6370 0.6320 ;
      RECT 5.6000 1.1790 6.3090 1.2290 ;
      RECT 5.5990 0.4500 5.6490 0.5630 ;
      RECT 5.5990 0.2970 5.6490 0.4000 ;
      RECT 5.6000 1.2290 5.6500 1.3530 ;
      RECT 5.1470 0.1880 5.7410 0.2380 ;
      RECT 5.1470 0.2380 5.1970 0.2880 ;
      RECT 4.5060 0.2880 5.1970 0.3380 ;
      RECT 4.1190 0.4550 4.1690 0.6130 ;
      RECT 3.6830 0.6130 4.1690 0.6630 ;
      RECT 4.5060 0.3380 4.5560 0.4050 ;
      RECT 4.1190 0.4050 4.5560 0.4550 ;
      RECT 6.9910 0.6130 7.4130 0.6630 ;
      RECT 6.3590 0.8090 6.4090 1.3010 ;
      RECT 6.3590 0.5500 6.4090 0.7590 ;
      RECT 6.1310 0.5000 6.4090 0.5500 ;
      RECT 6.1310 0.5500 6.1810 0.6790 ;
      RECT 6.6630 0.8090 6.7130 1.3010 ;
      RECT 6.9910 0.6630 7.0410 0.7590 ;
      RECT 6.3590 0.7590 7.0410 0.8090 ;
      RECT 3.0150 0.8130 3.1050 0.8630 ;
      RECT 3.0550 0.4620 3.1050 0.8130 ;
      RECT 3.0150 0.8630 3.0650 1.0830 ;
      RECT 2.9990 0.4120 3.1050 0.4620 ;
      RECT 2.2550 1.0830 3.0650 1.1330 ;
      RECT 3.0150 1.1330 3.0650 1.3540 ;
      RECT 2.2550 0.7520 2.3050 1.0830 ;
      RECT 2.2550 0.7020 2.3450 0.7520 ;
      RECT 2.2950 0.5510 2.3450 0.7020 ;
      RECT 2.2550 0.5010 2.3450 0.5510 ;
      RECT 2.2550 0.4070 2.3050 0.5010 ;
      RECT 2.4070 0.6130 2.8530 0.6630 ;
      RECT 2.4070 0.6630 2.4570 1.0040 ;
      RECT 2.4070 0.4130 2.4570 0.6130 ;
      RECT 6.4350 0.1380 6.4850 0.1700 ;
      RECT 3.5020 0.0880 6.4850 0.1380 ;
      RECT 8.3190 0.8200 8.8670 0.8700 ;
      RECT 1.6500 0.7020 1.9410 0.7280 ;
      RECT 1.6870 0.6780 1.9410 0.7020 ;
      RECT 1.3430 0.4600 1.3930 0.5020 ;
      RECT 1.0230 0.4100 1.3930 0.4600 ;
      RECT 1.0230 1.0200 1.7000 1.0700 ;
      RECT 1.6500 0.7520 1.7000 1.0200 ;
      RECT 1.6500 0.7280 1.7370 0.7520 ;
      RECT 1.6870 0.5520 1.7370 0.6780 ;
      RECT 1.3430 0.5020 1.7370 0.5520 ;
      RECT 0.8870 0.3100 1.5450 0.3600 ;
      RECT 1.4950 0.3600 1.5450 0.3920 ;
      RECT 0.8870 0.3600 0.9370 0.3920 ;
      RECT 5.6590 0.8660 5.8080 0.9160 ;
      RECT 5.7580 0.9160 5.8080 0.9670 ;
      RECT 5.7580 0.9670 5.8930 1.0170 ;
      RECT 1.9910 0.6280 2.2450 0.6520 ;
      RECT 1.9520 0.6020 2.2450 0.6280 ;
      RECT 1.9910 0.6520 2.0410 0.7780 ;
      RECT 1.9520 0.5780 2.0410 0.6020 ;
      RECT 1.9520 0.7780 2.0410 0.8280 ;
      RECT 1.9520 0.3190 2.0020 0.5780 ;
      RECT 1.9520 0.8280 2.0020 1.0760 ;
      RECT 8.6230 0.7090 9.1610 0.7590 ;
      RECT 4.6710 0.4880 5.2320 0.5110 ;
      RECT 4.6710 0.5110 5.2330 0.5380 ;
      RECT 5.1830 0.5380 5.2330 1.0200 ;
      RECT 4.6870 1.0200 5.2330 1.0700 ;
      RECT 4.4230 0.7880 4.4730 1.1200 ;
      RECT 3.3740 0.7380 4.4750 0.7880 ;
      RECT 4.2310 0.5050 4.2810 0.7380 ;
      RECT 4.6870 1.0700 4.7370 1.1200 ;
      RECT 3.9110 1.1200 4.7370 1.1700 ;
      RECT 5.2010 1.5200 8.3250 1.5700 ;
      RECT 9.2470 0.6770 9.2970 0.7680 ;
      RECT 9.2070 0.4270 9.2970 0.4620 ;
      RECT 9.2470 0.1260 9.2970 0.4270 ;
      RECT 9.2070 0.6270 9.2970 0.6770 ;
      RECT 9.2070 0.5120 9.2570 0.6270 ;
      RECT 9.0030 0.4770 9.2570 0.5120 ;
      RECT 9.0030 0.4620 9.2970 0.4770 ;
      RECT 4.4430 1.5200 5.1330 1.5700 ;
      RECT 4.8980 0.6130 5.1330 0.6630 ;
      RECT 5.4470 0.8670 5.5890 0.9170 ;
      RECT 5.4470 0.6630 5.4970 0.8670 ;
      RECT 5.4470 0.6130 5.8930 0.6630 ;
      RECT 4.5350 0.9200 4.9650 0.9700 ;
      RECT 4.9150 0.8310 4.9650 0.9200 ;
      RECT 4.5350 0.9700 4.5850 1.0340 ;
      RECT 4.5350 0.5050 4.5850 0.9200 ;
      RECT 4.2910 1.4200 5.5970 1.4700 ;
      RECT 3.3030 1.1900 3.6890 1.2400 ;
      RECT 5.8800 1.2790 6.2730 1.3290 ;
      RECT 2.9220 0.0940 3.3150 0.1440 ;
      RECT 3.2270 1.3890 3.7650 1.4390 ;
      RECT 7.3310 1.2390 8.6290 1.2890 ;
      RECT 7.9390 0.5270 8.5370 0.5770 ;
      RECT 8.4870 0.5770 8.5370 0.7700 ;
      RECT 8.4870 0.3480 8.5370 0.5270 ;
      RECT 8.1830 0.5770 8.2330 0.8800 ;
      RECT 8.1830 0.1260 8.2330 0.5270 ;
      RECT 8.6230 0.1320 8.8570 0.1820 ;
      RECT 7.8790 1.0970 8.3280 1.1470 ;
      RECT 7.8790 0.6770 7.9290 1.0970 ;
      RECT 7.8390 0.6270 7.9290 0.6770 ;
      RECT 7.8390 0.4770 7.8890 0.6270 ;
      RECT 7.8390 0.4270 7.9290 0.4770 ;
      RECT 7.8790 0.1260 7.9290 0.4270 ;
      RECT 2.6190 1.5240 3.9170 1.5740 ;
      RECT 0.7190 0.5100 1.2570 0.5600 ;
      RECT 1.1750 1.1330 1.5610 1.1830 ;
      RECT 0.7190 0.9410 0.9530 0.9910 ;
      RECT 8.8510 1.0970 9.3890 1.1470 ;
      RECT 8.3190 0.2480 9.1610 0.2980 ;
      RECT 2.8630 0.7130 2.9890 0.7630 ;
      RECT 2.8630 0.7630 2.9130 1.0330 ;
      RECT 2.9390 0.5630 2.9890 0.7130 ;
      RECT 2.8470 0.5130 2.9890 0.5630 ;
      RECT 4.8230 0.3880 5.4970 0.4380 ;
      RECT 5.4470 0.4380 5.4970 0.5630 ;
      RECT 5.4470 0.2970 5.4970 0.3880 ;
    LAYER PO ;
      RECT 9.4850 0.0660 9.5150 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 5.8370 0.0660 5.8670 0.6910 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 3.1010 0.8400 3.1310 1.6060 ;
      RECT 5.8370 0.9390 5.8670 1.6060 ;
      RECT 5.5330 0.0660 5.5630 0.6370 ;
      RECT 3.1010 0.0660 3.1310 0.6370 ;
      RECT 9.3330 0.0660 9.3630 1.6060 ;
      RECT 3.7090 0.0660 3.7390 0.6910 ;
      RECT 5.0770 0.0660 5.1070 0.6910 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 9.6370 0.0660 9.6670 1.6060 ;
      RECT 4.7730 0.8920 4.8030 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 5.5330 0.8390 5.5630 1.6060 ;
      RECT 9.7890 0.0660 9.8190 1.6060 ;
      RECT 10.2450 0.0660 10.2750 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 9.9410 0.0660 9.9710 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 10.0930 0.0660 10.1230 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 4.7730 0.0660 4.8030 0.6910 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 3.7090 0.9390 3.7390 1.6060 ;
      RECT 7.3570 0.0670 7.3870 1.6050 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 5.0770 0.8390 5.1070 1.6060 ;
    LAYER NWELL ;
      RECT 7.7120 0.4910 9.7230 1.0830 ;
      RECT -0.1150 1.5430 10.4580 1.7730 ;
      RECT -0.1150 0.6790 7.2500 1.5430 ;
      RECT 10.1830 0.6790 10.4580 1.5430 ;
  END
END RSDFFNSRASX1_LVT

MACRO RSDFFNSRASX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.64 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3770 1.4650 2.5490 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 10.6400 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 1.6470 1.1310 1.6970 1.6420 ;
        RECT 2.1030 1.1310 2.1530 1.6420 ;
        RECT 1.7990 1.1310 1.8490 1.6420 ;
        RECT 2.2550 1.2940 2.3050 1.6420 ;
        RECT 3.9670 1.2700 4.0170 1.6420 ;
        RECT 8.6790 1.4540 8.7290 1.6420 ;
        RECT 2.2550 1.2440 2.7770 1.2940 ;
        RECT 3.7580 1.2200 5.0570 1.2700 ;
        RECT 5.7510 1.4040 8.7290 1.4540 ;
        RECT 5.7510 1.2790 5.8010 1.4040 ;
        RECT 6.8150 0.9130 6.8650 1.4040 ;
        RECT 7.1190 0.9610 7.1690 1.4040 ;
        RECT 6.5110 0.9530 6.5610 1.4040 ;
        RECT 7.4230 1.0530 7.4730 1.4040 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 10.6400 0.0300 ;
        RECT 2.1030 0.0300 2.1530 0.3070 ;
        RECT 1.6470 0.0300 1.6970 0.4050 ;
        RECT 0.5830 0.0300 0.6330 0.5120 ;
        RECT 0.4310 0.0300 0.4810 0.4340 ;
        RECT 1.7990 0.0300 1.8490 0.4050 ;
        RECT 7.4230 0.0300 7.4730 0.2210 ;
        RECT 6.8150 0.0300 6.8650 0.4090 ;
        RECT 7.1190 0.0300 7.1690 0.3200 ;
        RECT 8.3350 0.0300 8.3850 0.4260 ;
        RECT 9.7030 0.0300 9.7530 0.4260 ;
        RECT 9.2470 0.0300 9.2970 0.1980 ;
        RECT 6.6870 0.0300 6.7370 0.2880 ;
        RECT 2.1030 0.3070 3.9770 0.3570 ;
        RECT 5.7350 0.2880 6.7370 0.3380 ;
        RECT 3.7750 0.3570 3.8250 0.5570 ;
        RECT 2.5590 0.3570 2.6090 0.5570 ;
        RECT 2.7110 0.3570 2.7610 0.5570 ;
        RECT 3.9270 0.3570 3.9770 0.5330 ;
        RECT 2.1030 0.3570 2.1530 0.4050 ;
        RECT 3.9270 0.2380 3.9770 0.3070 ;
        RECT 3.9270 0.1880 5.0570 0.2380 ;
        RECT 4.3830 0.2380 4.4330 0.3490 ;
    END
  END VSS

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.9790 0.8570 6.1350 0.9750 ;
        RECT 5.9790 0.9750 6.0290 1.0790 ;
        RECT 5.4470 1.0790 6.0290 1.1290 ;
        RECT 5.4470 1.1290 5.4970 1.3200 ;
        RECT 4.1550 1.3200 5.4970 1.3700 ;
        RECT 4.1550 1.3700 4.2050 1.4550 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.9670 0.8330 7.8190 0.8830 ;
        RECT 6.9670 0.8830 7.0170 1.3190 ;
        RECT 7.7690 0.5110 7.8190 0.8330 ;
        RECT 7.6970 0.4520 7.8190 0.5110 ;
        RECT 6.9670 0.4020 7.8190 0.4520 ;
        RECT 6.9670 0.1490 7.0170 0.4020 ;
        RECT 7.6970 0.4010 7.8190 0.4020 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.8250 0.2490 9.9350 0.3590 ;
        RECT 9.8360 0.3590 9.8860 0.5270 ;
        RECT 9.6110 0.5270 9.8860 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.7630 0.5970 4.8130 0.7050 ;
        RECT 4.6570 0.7050 4.8130 0.7310 ;
        RECT 4.6570 0.7310 5.1170 0.7810 ;
        RECT 4.6570 0.7810 4.8130 0.8150 ;
        RECT 5.0670 0.7810 5.1170 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.2710 0.2710 7.9690 0.3210 ;
        RECT 7.8490 0.3210 7.9690 0.3590 ;
        RECT 7.8490 0.2490 7.9690 0.2710 ;
        RECT 7.2710 0.1490 7.3210 0.2710 ;
        RECT 7.9190 0.3590 7.9690 0.9330 ;
        RECT 7.2710 0.9330 7.9690 0.9830 ;
        RECT 7.2710 0.9830 7.3210 1.3270 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 8.3190 0.9490 9.9370 1.0090 ;
        RECT 9.8270 0.6900 9.9370 0.9490 ;
        RECT 9.7030 0.6270 9.7530 0.9490 ;
    END
  END VDDG

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2520 1.3330 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6780 0.7250 0.7280 ;
        RECT 0.4010 0.5510 0.5110 0.6780 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 1.1610 1.0110 1.3160 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D
  OBS
    LAYER M1 ;
      RECT 6.4350 0.1380 6.4850 0.1700 ;
      RECT 3.5470 0.0880 6.4850 0.1380 ;
      RECT 3.5470 0.1380 3.5970 0.1700 ;
      RECT 1.4520 0.6020 1.6370 0.6520 ;
      RECT 0.2050 0.8410 1.5020 0.8910 ;
      RECT 1.4520 0.6520 1.5020 0.8410 ;
      RECT 0.2050 0.5260 0.2550 0.8410 ;
      RECT 0.2790 0.8910 0.3290 1.2140 ;
      RECT 0.2050 0.4760 0.3290 0.5260 ;
      RECT 0.2790 0.3160 0.3290 0.4760 ;
      RECT 0.8870 0.3100 1.5450 0.3600 ;
      RECT 1.4950 0.3600 1.5450 0.3920 ;
      RECT 0.8870 0.3600 0.9370 0.3920 ;
      RECT 1.6870 0.6780 1.9410 0.7020 ;
      RECT 1.6500 0.7020 1.9410 0.7280 ;
      RECT 1.3430 0.4600 1.3930 0.5020 ;
      RECT 1.0230 0.4100 1.3930 0.4600 ;
      RECT 1.3430 0.5020 1.7370 0.5520 ;
      RECT 1.6870 0.5520 1.7370 0.6780 ;
      RECT 1.6500 0.7280 1.7370 0.7520 ;
      RECT 1.6500 0.7520 1.7000 1.0200 ;
      RECT 1.0230 1.0200 1.7000 1.0700 ;
      RECT 0.7190 0.5100 1.2570 0.5600 ;
      RECT 3.1670 0.8540 4.0690 0.9040 ;
      RECT 3.1670 0.4130 3.2170 0.5630 ;
      RECT 3.1670 0.5630 3.3690 0.6130 ;
      RECT 3.1670 0.6130 3.2170 0.8540 ;
      RECT 3.3190 0.4070 3.3690 0.5630 ;
      RECT 3.1670 0.9040 3.2170 1.0590 ;
      RECT 3.1670 1.0590 3.5370 1.1090 ;
      RECT 3.1670 1.1090 3.2170 1.3370 ;
      RECT 1.9910 0.6280 2.2450 0.6520 ;
      RECT 1.9520 0.6020 2.2450 0.6280 ;
      RECT 1.9910 0.6520 2.0410 0.7780 ;
      RECT 1.9520 0.5780 2.0410 0.6020 ;
      RECT 1.9520 0.7780 2.0410 0.8280 ;
      RECT 1.9520 0.3190 2.0020 0.5780 ;
      RECT 1.9520 0.8280 2.0020 1.0760 ;
      RECT 2.8470 0.5130 2.9890 0.5630 ;
      RECT 2.9390 0.5630 2.9890 0.7130 ;
      RECT 2.8630 0.7130 2.9890 0.7630 ;
      RECT 2.8630 0.7630 2.9130 1.0330 ;
      RECT 2.9990 0.4120 3.1050 0.4620 ;
      RECT 3.0550 0.4620 3.1050 0.8130 ;
      RECT 3.0150 0.8130 3.1050 0.8630 ;
      RECT 3.0150 0.8630 3.0650 1.0830 ;
      RECT 2.2550 1.0830 3.0650 1.1330 ;
      RECT 3.0150 1.1330 3.0650 1.3540 ;
      RECT 2.2550 0.7520 2.3050 1.0830 ;
      RECT 2.2550 0.7020 2.3450 0.7520 ;
      RECT 2.2950 0.5510 2.3450 0.7020 ;
      RECT 2.2550 0.5010 2.3450 0.5510 ;
      RECT 2.2550 0.4070 2.3050 0.5010 ;
      RECT 2.4070 0.6130 2.8530 0.6630 ;
      RECT 2.4070 0.6630 2.4570 1.0040 ;
      RECT 2.4070 0.4130 2.4570 0.6130 ;
      RECT 2.9220 0.0940 3.3150 0.1440 ;
      RECT 5.1470 0.1880 5.7410 0.2380 ;
      RECT 5.1470 0.2380 5.1970 0.2880 ;
      RECT 4.5060 0.2880 5.1970 0.3380 ;
      RECT 4.1190 0.4550 4.1690 0.6130 ;
      RECT 3.6830 0.6130 4.1690 0.6630 ;
      RECT 4.5060 0.3380 4.5560 0.4050 ;
      RECT 4.1190 0.4050 4.5560 0.4550 ;
      RECT 4.8230 0.3880 5.4970 0.4380 ;
      RECT 5.4470 0.4380 5.4970 0.5630 ;
      RECT 5.4470 0.2970 5.4970 0.3880 ;
      RECT 5.2950 0.9670 5.5130 1.0170 ;
      RECT 5.2950 0.4380 5.3450 0.9670 ;
      RECT 5.2950 1.0170 5.3450 1.1200 ;
      RECT 5.2950 1.1700 5.3450 1.2700 ;
      RECT 4.8230 1.1200 5.3450 1.1700 ;
      RECT 6.5690 0.6320 7.1090 0.6820 ;
      RECT 5.9430 0.4500 5.9930 0.7290 ;
      RECT 5.9430 0.7290 6.3090 0.7790 ;
      RECT 6.2590 0.7790 6.3090 1.1790 ;
      RECT 6.5870 0.4500 6.6370 0.6320 ;
      RECT 5.5990 0.4000 6.6370 0.4500 ;
      RECT 5.6000 1.1790 6.3090 1.2290 ;
      RECT 5.5990 0.4500 5.6490 0.5630 ;
      RECT 5.5990 0.2970 5.6490 0.4000 ;
      RECT 5.6000 1.2290 5.6500 1.3530 ;
      RECT 5.1830 0.5380 5.2330 1.0200 ;
      RECT 4.6710 0.5110 5.2330 0.5380 ;
      RECT 4.6870 1.0200 5.2330 1.0700 ;
      RECT 4.6710 0.4880 5.2320 0.5110 ;
      RECT 4.4230 0.7880 4.4730 1.1200 ;
      RECT 3.3740 0.7380 4.4750 0.7880 ;
      RECT 4.2310 0.5050 4.2810 0.7380 ;
      RECT 4.6870 1.0700 4.7370 1.1200 ;
      RECT 3.9110 1.1200 4.7370 1.1700 ;
      RECT 4.8980 0.6130 5.1330 0.6630 ;
      RECT 5.4470 0.6130 5.8930 0.6630 ;
      RECT 5.4470 0.6630 5.4970 0.8670 ;
      RECT 5.4470 0.8670 5.5890 0.9170 ;
      RECT 4.5350 0.9200 4.9650 0.9700 ;
      RECT 4.9150 0.8310 4.9650 0.9200 ;
      RECT 4.5350 0.9700 4.5850 1.0340 ;
      RECT 4.5350 0.5050 4.5850 0.9200 ;
      RECT 7.1790 0.6130 7.7170 0.6630 ;
      RECT 7.1790 0.6630 7.2290 0.7320 ;
      RECT 6.3590 0.7320 7.2290 0.7820 ;
      RECT 6.3590 0.7820 6.4090 1.3010 ;
      RECT 6.3590 0.5500 6.4090 0.7320 ;
      RECT 6.1310 0.5000 6.4090 0.5500 ;
      RECT 6.1310 0.5500 6.1810 0.6790 ;
      RECT 6.6630 0.7820 6.7130 1.3010 ;
      RECT 8.1830 1.0840 8.6320 1.1340 ;
      RECT 8.1830 0.6770 8.2330 1.0840 ;
      RECT 8.1430 0.6270 8.2330 0.6770 ;
      RECT 8.1430 0.4770 8.1930 0.6270 ;
      RECT 8.1430 0.4270 8.2330 0.4770 ;
      RECT 8.1830 0.1260 8.2330 0.4270 ;
      RECT 8.2430 0.5270 8.8410 0.5770 ;
      RECT 8.7910 0.5770 8.8410 0.7700 ;
      RECT 8.7910 0.3480 8.8410 0.5270 ;
      RECT 8.4870 0.5770 8.5370 0.8870 ;
      RECT 8.4870 0.1260 8.5370 0.5270 ;
      RECT 8.6230 0.2480 9.4650 0.2980 ;
      RECT 9.5510 0.6770 9.6010 0.7680 ;
      RECT 9.5110 0.4270 9.6010 0.4620 ;
      RECT 9.5510 0.1260 9.6010 0.4270 ;
      RECT 9.5110 0.6270 9.6010 0.6770 ;
      RECT 9.5110 0.5120 9.5610 0.6270 ;
      RECT 9.3070 0.4770 9.5610 0.5120 ;
      RECT 9.3070 0.4620 9.6010 0.4770 ;
      RECT 8.9270 0.1320 9.1610 0.1820 ;
      RECT 1.1750 1.1330 1.5610 1.1830 ;
      RECT 0.7190 0.9410 0.9530 0.9910 ;
      RECT 3.3030 1.1900 3.6890 1.2400 ;
      RECT 3.2270 1.3890 3.7650 1.4390 ;
      RECT 3.6830 0.9680 4.2630 1.0180 ;
      RECT 4.2130 0.9080 4.2630 0.9680 ;
      RECT 4.2130 0.8580 4.3730 0.9080 ;
      RECT 2.6190 1.5240 3.9170 1.5740 ;
      RECT 5.7580 0.9670 5.8930 1.0170 ;
      RECT 5.7580 0.9160 5.8080 0.9670 ;
      RECT 5.6590 0.8660 5.8080 0.9160 ;
      RECT 4.4430 1.5200 5.1330 1.5700 ;
      RECT 4.2910 1.4200 5.5970 1.4700 ;
      RECT 5.8800 1.2790 6.2730 1.3290 ;
      RECT 7.6350 1.2230 8.9330 1.2730 ;
      RECT 8.6230 0.8200 9.1710 0.8700 ;
      RECT 8.9270 0.7090 9.4650 0.7590 ;
      RECT 9.1550 1.0820 9.6930 1.1320 ;
      RECT 5.2010 1.5200 8.6290 1.5700 ;
    LAYER PO ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 3.7090 0.9390 3.7390 1.6060 ;
      RECT 7.6610 0.0670 7.6910 1.6050 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 9.3330 0.0660 9.3630 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 5.0770 0.8390 5.1070 1.6060 ;
      RECT 9.7890 0.0660 9.8190 1.6060 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 9.4850 0.0660 9.5150 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 5.8370 0.0660 5.8670 0.6910 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 3.1010 0.8400 3.1310 1.6060 ;
      RECT 5.8370 0.9390 5.8670 1.6060 ;
      RECT 5.5330 0.0660 5.5630 0.6370 ;
      RECT 3.7090 0.0660 3.7390 0.6910 ;
      RECT 3.1010 0.0660 3.1310 0.6370 ;
      RECT 9.6370 0.0660 9.6670 1.6060 ;
      RECT 5.0770 0.0660 5.1070 0.6910 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 9.9410 0.0660 9.9710 1.6060 ;
      RECT 4.7730 0.8920 4.8030 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 5.5330 0.8390 5.5630 1.6060 ;
      RECT 10.0930 0.0660 10.1230 1.6060 ;
      RECT 10.5490 0.0660 10.5790 1.6060 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 10.2450 0.0660 10.2750 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 10.3970 0.0660 10.4270 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 4.7730 0.0660 4.8030 0.6910 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
    LAYER NWELL ;
      RECT 8.0160 0.4910 10.0270 1.0830 ;
      RECT -0.1150 1.5430 10.7620 1.7730 ;
      RECT -0.1150 0.6790 7.5540 1.5430 ;
      RECT 10.4870 0.6790 10.7620 1.5430 ;
  END
END RSDFFNSRASX2_LVT

MACRO RSDFFNSRX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.728 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 9.7280 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 2.1030 1.1310 2.1530 1.6420 ;
        RECT 1.7990 1.1310 1.8490 1.6420 ;
        RECT 1.6470 1.1310 1.6970 1.6420 ;
        RECT 2.2550 1.2940 2.3050 1.6420 ;
        RECT 3.8150 1.2700 3.8650 1.6420 ;
        RECT 7.7670 1.4540 7.8170 1.6420 ;
        RECT 2.2550 1.2440 2.7770 1.2940 ;
        RECT 3.6070 1.2200 4.7530 1.2700 ;
        RECT 5.4470 1.4040 7.8170 1.4540 ;
        RECT 5.4470 1.2790 5.4970 1.4040 ;
        RECT 6.3590 0.9590 6.4090 1.4040 ;
        RECT 5.9030 0.9530 5.9530 1.4040 ;
    END
  END VDD

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.2070 0.4010 6.9070 0.4510 ;
        RECT 6.2070 0.1570 6.2570 0.4010 ;
        RECT 6.7850 0.4510 6.9070 0.5380 ;
        RECT 6.8570 0.5380 6.9070 0.8590 ;
        RECT 6.2070 0.8590 6.9070 0.9090 ;
        RECT 6.2070 0.9090 6.2570 1.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.5110 0.9690 7.0450 1.0190 ;
        RECT 6.9950 0.3510 7.0450 0.9690 ;
        RECT 6.5110 1.0190 6.7430 1.1290 ;
        RECT 6.4950 0.3010 7.0450 0.3510 ;
        RECT 6.5110 1.1290 6.5610 1.3270 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3770 1.4650 2.5490 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 9.7280 0.0300 ;
        RECT 2.1030 0.0300 2.1530 0.2570 ;
        RECT 8.7910 0.0300 8.8410 0.4260 ;
        RECT 1.6470 0.0300 1.6970 0.4050 ;
        RECT 6.3590 0.0300 6.4090 0.2410 ;
        RECT 1.7990 0.0300 1.8490 0.4050 ;
        RECT 7.4230 0.0300 7.4730 0.4260 ;
        RECT 0.5830 0.0300 0.6330 0.5120 ;
        RECT 0.4310 0.0300 0.4810 0.4340 ;
        RECT 8.3350 0.0300 8.3850 0.1980 ;
        RECT 6.0790 0.0300 6.1290 0.2830 ;
        RECT 2.1030 0.2570 3.8250 0.3070 ;
        RECT 5.4310 0.2830 6.1290 0.3330 ;
        RECT 2.5590 0.3070 2.6090 0.5570 ;
        RECT 2.7110 0.3070 2.7610 0.5570 ;
        RECT 2.1030 0.3070 2.1530 0.4050 ;
        RECT 3.7750 0.2340 3.8250 0.2570 ;
        RECT 3.7750 0.1840 4.7530 0.2340 ;
        RECT 4.0790 0.2340 4.1290 0.3490 ;
    END
  END VSS

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.9130 0.2490 9.0230 0.3590 ;
        RECT 8.9240 0.3590 8.9740 0.5170 ;
        RECT 8.6990 0.5170 8.9740 0.5670 ;
        RECT 8.9240 0.5670 8.9740 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.3530 0.7050 4.5090 0.7310 ;
        RECT 4.3530 0.7310 4.8130 0.7810 ;
        RECT 4.4590 0.5970 4.5090 0.7050 ;
        RECT 4.3530 0.7810 4.5090 0.8150 ;
        RECT 4.7630 0.7810 4.8130 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 7.4070 0.9510 9.0250 1.0110 ;
        RECT 8.9150 0.6900 9.0250 0.9510 ;
        RECT 8.7910 0.6270 8.8410 0.9510 ;
    END
  END VDDG

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2520 1.3330 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6780 0.7250 0.7280 ;
        RECT 0.4010 0.5510 0.5110 0.6780 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 1.1610 1.0110 1.3160 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D
  OBS
    LAYER M1 ;
      RECT 5.2960 1.2290 5.3460 1.3530 ;
      RECT 1.6500 0.7020 1.9410 0.7280 ;
      RECT 1.6870 0.6780 1.9410 0.7020 ;
      RECT 1.3430 0.4600 1.3930 0.5020 ;
      RECT 1.0230 0.4100 1.3930 0.4600 ;
      RECT 1.0230 1.0200 1.7000 1.0700 ;
      RECT 1.6500 0.7520 1.7000 1.0200 ;
      RECT 1.6500 0.7280 1.7370 0.7520 ;
      RECT 1.6870 0.5520 1.7370 0.6780 ;
      RECT 1.3430 0.5020 1.7370 0.5520 ;
      RECT 0.8870 0.3100 1.5450 0.3600 ;
      RECT 1.4950 0.3600 1.5450 0.3920 ;
      RECT 0.8870 0.3600 0.9370 0.3920 ;
      RECT 5.3550 0.8660 5.5040 0.9160 ;
      RECT 5.4540 0.9160 5.5040 0.9670 ;
      RECT 5.4540 0.9670 5.5890 1.0170 ;
      RECT 6.3830 0.6130 6.8050 0.6630 ;
      RECT 6.0550 0.8090 6.1050 1.3010 ;
      RECT 5.8270 0.5670 5.8770 0.7590 ;
      RECT 5.8260 0.5170 5.9690 0.5670 ;
      RECT 6.3830 0.6630 6.4330 0.7590 ;
      RECT 5.8260 0.7590 6.4330 0.8090 ;
      RECT 1.9910 0.6280 2.2450 0.6520 ;
      RECT 1.9520 0.6020 2.2450 0.6280 ;
      RECT 1.9910 0.6520 2.0410 0.7780 ;
      RECT 1.9520 0.5780 2.0410 0.6020 ;
      RECT 1.9520 0.7780 2.0410 0.8280 ;
      RECT 1.9520 0.3190 2.0020 0.5780 ;
      RECT 1.9520 0.8280 2.0020 1.0760 ;
      RECT 2.2550 1.0830 3.0650 1.1330 ;
      RECT 3.0150 1.1330 3.0650 1.3540 ;
      RECT 3.0150 0.8630 3.0650 1.0830 ;
      RECT 3.0150 0.8130 3.1050 0.8630 ;
      RECT 3.0550 0.4620 3.1050 0.8130 ;
      RECT 2.9990 0.4120 3.1050 0.4620 ;
      RECT 2.2550 0.7520 2.3050 1.0830 ;
      RECT 2.2550 0.7020 2.3450 0.7520 ;
      RECT 2.2950 0.5510 2.3450 0.7020 ;
      RECT 2.2550 0.5010 2.3450 0.5510 ;
      RECT 2.2550 0.4070 2.3050 0.5010 ;
      RECT 8.0150 0.7090 8.5530 0.7590 ;
      RECT 3.2270 1.4240 3.6130 1.4740 ;
      RECT 3.1670 0.8540 3.9170 0.9040 ;
      RECT 3.1670 0.4840 3.2170 0.8540 ;
      RECT 3.1670 0.9040 3.2170 1.0990 ;
      RECT 3.1670 0.4340 3.3850 0.4840 ;
      RECT 3.1670 1.0990 3.3850 1.1490 ;
      RECT 3.1670 0.4080 3.2170 0.4340 ;
      RECT 3.1670 1.1490 3.2170 1.3370 ;
      RECT 2.4070 0.6130 2.8530 0.6630 ;
      RECT 2.4070 0.6630 2.4570 1.0040 ;
      RECT 2.4070 0.4130 2.4570 0.6130 ;
      RECT 4.8790 0.5340 4.9290 1.0200 ;
      RECT 4.3670 0.5070 4.9290 0.5340 ;
      RECT 4.3830 1.0200 4.9290 1.0700 ;
      RECT 4.3670 0.4840 4.9280 0.5070 ;
      RECT 4.1190 0.7880 4.1690 1.1200 ;
      RECT 3.3730 0.7380 4.1710 0.7880 ;
      RECT 3.9270 0.5050 3.9770 0.7380 ;
      RECT 4.3830 1.0700 4.4330 1.1200 ;
      RECT 3.7590 1.1200 4.4330 1.1700 ;
      RECT 8.5990 0.6270 8.6890 0.6770 ;
      RECT 8.6390 0.6770 8.6890 0.7680 ;
      RECT 8.5990 0.4530 8.6490 0.4620 ;
      RECT 8.5990 0.4030 8.6890 0.4530 ;
      RECT 8.6390 0.1260 8.6890 0.4030 ;
      RECT 8.5990 0.5120 8.6490 0.6270 ;
      RECT 8.3950 0.4620 8.6490 0.5120 ;
      RECT 4.1390 1.5200 4.8290 1.5700 ;
      RECT 4.5940 0.6130 4.8290 0.6630 ;
      RECT 5.1430 0.8670 5.2850 0.9170 ;
      RECT 5.1430 0.6630 5.1930 0.8670 ;
      RECT 5.1430 0.6130 5.5890 0.6630 ;
      RECT 4.8430 0.1780 5.4370 0.2280 ;
      RECT 4.8430 0.2280 4.8930 0.2840 ;
      RECT 4.2020 0.2840 4.8930 0.3340 ;
      RECT 3.5470 0.5240 3.5970 0.6130 ;
      RECT 3.7820 0.4550 3.8320 0.6130 ;
      RECT 3.5470 0.6130 3.8320 0.6630 ;
      RECT 4.2020 0.3340 4.2520 0.4050 ;
      RECT 3.7820 0.4050 4.2520 0.4550 ;
      RECT 4.2310 0.9200 4.6610 0.9700 ;
      RECT 4.6110 0.8310 4.6610 0.9200 ;
      RECT 4.2310 0.9700 4.2810 1.0340 ;
      RECT 4.2310 0.5050 4.2810 0.9200 ;
      RECT 3.9870 1.4200 5.2930 1.4700 ;
      RECT 6.7230 1.2190 8.0210 1.2690 ;
      RECT 2.9220 0.0940 3.3150 0.1440 ;
      RECT 7.7110 0.8200 8.2590 0.8700 ;
      RECT 8.0150 0.1320 8.2490 0.1820 ;
      RECT 7.2710 1.0780 7.7200 1.1280 ;
      RECT 7.2710 0.6770 7.3210 1.0780 ;
      RECT 7.2310 0.6270 7.3210 0.6770 ;
      RECT 7.2310 0.4770 7.2810 0.6270 ;
      RECT 7.2310 0.4270 7.3210 0.4770 ;
      RECT 7.2710 0.1260 7.3210 0.4270 ;
      RECT 2.6190 1.5240 3.7650 1.5740 ;
      RECT 7.3310 0.5270 7.9290 0.5770 ;
      RECT 7.5750 0.5770 7.6250 0.8870 ;
      RECT 7.5750 0.1260 7.6250 0.5270 ;
      RECT 7.8790 0.5770 7.9290 0.7700 ;
      RECT 7.8790 0.3480 7.9290 0.5270 ;
      RECT 5.6590 0.0880 5.8930 0.1380 ;
      RECT 0.7190 0.5100 1.2570 0.5600 ;
      RECT 1.1750 1.1330 1.5610 1.1830 ;
      RECT 0.7190 0.9410 0.9530 0.9910 ;
      RECT 8.2430 1.1060 8.7810 1.1560 ;
      RECT 7.7110 0.2480 8.5530 0.2980 ;
      RECT 4.8970 1.5200 7.7170 1.5700 ;
      RECT 2.8630 0.7130 2.9890 0.7630 ;
      RECT 2.8630 0.7630 2.9130 1.0330 ;
      RECT 2.9390 0.5630 2.9890 0.7130 ;
      RECT 2.8470 0.5130 2.9890 0.5630 ;
      RECT 4.5190 0.3840 5.1930 0.4340 ;
      RECT 5.1430 0.4340 5.1930 0.5630 ;
      RECT 5.1430 0.2970 5.1930 0.3840 ;
      RECT 4.9910 0.4340 5.0410 0.9670 ;
      RECT 4.9910 0.9670 5.2090 1.0170 ;
      RECT 4.9910 1.0170 5.0410 1.1200 ;
      RECT 4.9910 1.1700 5.0410 1.2700 ;
      RECT 4.5190 1.1200 5.0410 1.1700 ;
      RECT 3.5270 0.9680 4.0390 1.0180 ;
      RECT 3.9860 0.9080 4.0360 0.9680 ;
      RECT 3.9860 0.8580 4.0690 0.9080 ;
      RECT 1.4520 0.6020 1.6370 0.6520 ;
      RECT 0.2050 0.8410 1.5020 0.8910 ;
      RECT 1.4520 0.6520 1.5020 0.8410 ;
      RECT 0.2050 0.5260 0.2550 0.8410 ;
      RECT 0.2790 0.8910 0.3290 1.2140 ;
      RECT 0.2050 0.4760 0.3290 0.5260 ;
      RECT 0.2790 0.3160 0.3290 0.4760 ;
      RECT 5.9630 0.6320 6.3330 0.6820 ;
      RECT 6.2830 0.5970 6.3330 0.6320 ;
      RECT 5.6600 0.4500 5.7100 1.1790 ;
      RECT 5.2960 1.1790 5.8170 1.2290 ;
      RECT 6.0890 0.4500 6.1390 0.6320 ;
      RECT 5.2950 0.4000 6.1390 0.4500 ;
      RECT 5.2950 0.4500 5.3450 0.5630 ;
      RECT 5.2950 0.2970 5.3450 0.4000 ;
    LAYER PO ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.7090 0.0660 3.7390 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 3.1010 0.8400 3.1310 1.6060 ;
      RECT 5.5330 0.9390 5.5630 1.6060 ;
      RECT 5.2290 0.0660 5.2590 0.6370 ;
      RECT 3.1010 0.0660 3.1310 0.6370 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 4.7730 0.0660 4.8030 0.6910 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 4.4690 0.8920 4.4990 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 5.2290 0.8390 5.2590 1.6060 ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 9.6370 0.0660 9.6670 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 9.3330 0.0660 9.3630 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 9.4850 0.0660 9.5150 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 3.5570 0.0680 3.5870 0.6180 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 4.4690 0.0660 4.4990 0.6910 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 6.7490 0.0670 6.7790 1.6050 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 4.7730 0.8390 4.8030 1.6060 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 3.5570 0.7300 3.5870 1.6060 ;
      RECT 5.5330 0.0660 5.5630 0.6910 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
    LAYER NWELL ;
      RECT 7.1040 0.4910 9.1150 1.0830 ;
      RECT -0.1150 1.5430 9.8500 1.7730 ;
      RECT -0.1150 0.6790 6.6420 1.5430 ;
      RECT 9.5750 0.6790 9.8500 1.5430 ;
  END
END RSDFFNSRX1_LVT

MACRO RSDFFNSRX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.032 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 10.0320 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 2.1030 1.1310 2.1530 1.6420 ;
        RECT 1.7990 1.1310 1.8490 1.6420 ;
        RECT 1.6470 1.1310 1.6970 1.6420 ;
        RECT 8.0710 1.4540 8.1210 1.6420 ;
        RECT 2.2550 1.2940 2.3050 1.6420 ;
        RECT 3.8150 1.2700 3.8650 1.6420 ;
        RECT 5.4470 1.4040 8.1210 1.4540 ;
        RECT 2.2550 1.2440 2.7770 1.2940 ;
        RECT 3.6070 1.2200 4.7530 1.2700 ;
        RECT 5.4470 1.2790 5.4970 1.4040 ;
        RECT 5.9030 0.9530 5.9530 1.4040 ;
        RECT 6.2070 0.9130 6.2570 1.4040 ;
        RECT 6.5110 0.9610 6.5610 1.4040 ;
        RECT 6.8150 1.0530 6.8650 1.4040 ;
    END
  END VDD

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3770 1.4650 2.5490 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 10.0320 0.0300 ;
        RECT 2.1030 0.0300 2.1530 0.2570 ;
        RECT 6.8150 0.0300 6.8650 0.2210 ;
        RECT 9.0950 0.0300 9.1450 0.4260 ;
        RECT 1.6470 0.0300 1.6970 0.4050 ;
        RECT 6.5110 0.0300 6.5610 0.3200 ;
        RECT 6.2070 0.0300 6.2570 0.4090 ;
        RECT 1.7990 0.0300 1.8490 0.4050 ;
        RECT 7.7270 0.0300 7.7770 0.4260 ;
        RECT 0.5830 0.0300 0.6330 0.5120 ;
        RECT 0.4310 0.0300 0.4810 0.4340 ;
        RECT 8.6390 0.0300 8.6890 0.1980 ;
        RECT 6.0790 0.0300 6.1290 0.2830 ;
        RECT 2.1030 0.2570 3.8250 0.3070 ;
        RECT 5.4310 0.2830 6.1290 0.3330 ;
        RECT 2.5590 0.3070 2.6090 0.5570 ;
        RECT 2.7110 0.3070 2.7610 0.5570 ;
        RECT 2.1030 0.3070 2.1530 0.4050 ;
        RECT 3.7750 0.2340 3.8250 0.2570 ;
        RECT 3.7750 0.1840 4.7530 0.2340 ;
        RECT 4.0790 0.2340 4.1290 0.3490 ;
    END
  END VSS

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.2190 0.2490 9.3290 0.3590 ;
        RECT 9.2280 0.3590 9.2780 0.5270 ;
        RECT 9.0030 0.5270 9.2780 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.3530 0.7160 4.5090 0.7310 ;
        RECT 4.3530 0.7310 4.8130 0.7810 ;
        RECT 4.4590 0.5970 4.5090 0.7160 ;
        RECT 4.3530 0.7810 4.5090 0.8150 ;
        RECT 4.7630 0.7810 4.8130 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.6630 0.1490 6.7130 0.2710 ;
        RECT 6.6630 0.2710 7.3610 0.3210 ;
        RECT 7.2400 0.3210 7.3610 0.3600 ;
        RECT 7.2400 0.2500 7.3610 0.2710 ;
        RECT 7.3110 0.3600 7.3610 0.9330 ;
        RECT 6.6630 0.9330 7.3610 0.9830 ;
        RECT 6.6630 0.9830 6.7130 1.3270 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 7.7110 0.9470 9.3290 0.9970 ;
        RECT 9.2190 0.6900 9.3290 0.9470 ;
        RECT 9.0950 0.6270 9.1450 0.9470 ;
    END
  END VDDG

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.3590 0.8330 7.2110 0.8830 ;
        RECT 6.3590 0.8830 6.4090 1.3190 ;
        RECT 7.1610 0.5120 7.2110 0.8330 ;
        RECT 7.0890 0.4520 7.2110 0.5120 ;
        RECT 6.3590 0.4020 7.2110 0.4520 ;
        RECT 6.3590 0.1490 6.4090 0.4020 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2520 1.3330 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6780 0.7250 0.7280 ;
        RECT 0.4010 0.5510 0.5110 0.6780 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 1.1610 1.0110 1.3160 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D
  OBS
    LAYER M1 ;
      RECT 6.0890 0.4500 6.1390 0.6320 ;
      RECT 5.2950 0.4000 6.1390 0.4500 ;
      RECT 2.9990 0.4120 3.1050 0.4620 ;
      RECT 3.0550 0.4620 3.1050 0.8130 ;
      RECT 3.0150 0.8130 3.1050 0.8630 ;
      RECT 3.0150 0.8630 3.0650 1.0830 ;
      RECT 2.2550 1.0830 3.0650 1.1330 ;
      RECT 3.0150 1.1330 3.0650 1.3540 ;
      RECT 2.2550 0.7520 2.3050 1.0830 ;
      RECT 2.2550 0.7020 2.3450 0.7520 ;
      RECT 2.2950 0.5510 2.3450 0.7020 ;
      RECT 2.2550 0.5010 2.3450 0.5510 ;
      RECT 2.2550 0.4070 2.3050 0.5010 ;
      RECT 2.4070 0.6130 2.8530 0.6630 ;
      RECT 2.4070 0.6630 2.4570 1.0040 ;
      RECT 2.4070 0.4130 2.4570 0.6130 ;
      RECT 2.9220 0.0940 3.3150 0.1440 ;
      RECT 8.0150 0.8200 8.5630 0.8700 ;
      RECT 3.1670 0.8540 3.9170 0.9040 ;
      RECT 3.1670 0.4840 3.2170 0.8540 ;
      RECT 3.1670 0.9040 3.2170 1.0990 ;
      RECT 3.1670 0.4340 3.3850 0.4840 ;
      RECT 3.1670 1.0990 3.3850 1.1490 ;
      RECT 3.1670 0.4080 3.2170 0.4340 ;
      RECT 3.1670 1.1490 3.2170 1.3370 ;
      RECT 1.6500 0.7020 1.9410 0.7280 ;
      RECT 1.6870 0.6780 1.9410 0.7020 ;
      RECT 1.3430 0.4600 1.3930 0.5020 ;
      RECT 1.0230 0.4100 1.3930 0.4600 ;
      RECT 1.0230 1.0200 1.7000 1.0700 ;
      RECT 1.6500 0.7520 1.7000 1.0200 ;
      RECT 1.6500 0.7280 1.7370 0.7520 ;
      RECT 1.6870 0.5520 1.7370 0.6780 ;
      RECT 1.3430 0.5020 1.7370 0.5520 ;
      RECT 0.8870 0.3100 1.5450 0.3600 ;
      RECT 1.4950 0.3600 1.5450 0.3920 ;
      RECT 0.8870 0.3600 0.9370 0.3920 ;
      RECT 5.3550 0.8660 5.5040 0.9160 ;
      RECT 5.4540 0.9160 5.5040 0.9670 ;
      RECT 5.4540 0.9670 5.5890 1.0170 ;
      RECT 6.5620 0.6130 7.1090 0.6630 ;
      RECT 5.8270 0.7820 5.8770 0.8090 ;
      RECT 5.8270 0.5670 5.8770 0.7320 ;
      RECT 6.0550 0.7820 6.1050 1.3010 ;
      RECT 5.8260 0.5170 5.9690 0.5670 ;
      RECT 6.5620 0.6630 6.6120 0.7320 ;
      RECT 5.8260 0.7320 6.6120 0.7820 ;
      RECT 1.9910 0.6280 2.2450 0.6520 ;
      RECT 1.9520 0.6020 2.2450 0.6280 ;
      RECT 1.9910 0.6520 2.0410 0.7780 ;
      RECT 1.9520 0.5780 2.0410 0.6020 ;
      RECT 1.9520 0.7780 2.0410 0.8280 ;
      RECT 1.9520 0.3190 2.0020 0.5780 ;
      RECT 1.9520 0.8280 2.0020 1.0760 ;
      RECT 8.3190 0.7090 8.8570 0.7590 ;
      RECT 3.2270 1.4240 3.6130 1.4740 ;
      RECT 8.5470 1.0570 9.0850 1.1070 ;
      RECT 8.0150 0.2480 8.8570 0.2980 ;
      RECT 4.8790 0.5340 4.9290 1.0200 ;
      RECT 4.3670 0.5070 4.9290 0.5340 ;
      RECT 4.3830 1.0200 4.9290 1.0700 ;
      RECT 4.3670 0.4840 4.9280 0.5070 ;
      RECT 4.1190 0.7880 4.1690 1.1200 ;
      RECT 3.3730 0.7380 4.1710 0.7880 ;
      RECT 3.9270 0.5050 3.9770 0.7380 ;
      RECT 4.3830 1.0700 4.4330 1.1200 ;
      RECT 3.7590 1.1200 4.4330 1.1700 ;
      RECT 4.8970 1.5200 8.0210 1.5700 ;
      RECT 8.9430 0.6770 8.9930 0.7680 ;
      RECT 8.9030 0.4270 8.9930 0.4620 ;
      RECT 8.9430 0.1260 8.9930 0.4270 ;
      RECT 8.9030 0.6270 8.9930 0.6770 ;
      RECT 8.9030 0.5120 8.9530 0.6270 ;
      RECT 8.6990 0.4770 8.9530 0.5120 ;
      RECT 8.6990 0.4620 8.9930 0.4770 ;
      RECT 4.1390 1.5200 4.8290 1.5700 ;
      RECT 4.5940 0.6130 4.8290 0.6630 ;
      RECT 5.1430 0.8670 5.2850 0.9170 ;
      RECT 5.1430 0.6630 5.1930 0.8670 ;
      RECT 5.1430 0.6130 5.5890 0.6630 ;
      RECT 4.8430 0.1780 5.4370 0.2280 ;
      RECT 4.8430 0.2280 4.8930 0.2840 ;
      RECT 4.2020 0.2840 4.8930 0.3340 ;
      RECT 3.5470 0.5240 3.5970 0.6130 ;
      RECT 3.7820 0.4550 3.8320 0.6130 ;
      RECT 3.5470 0.6130 3.8320 0.6630 ;
      RECT 4.2020 0.3340 4.2520 0.4050 ;
      RECT 3.7820 0.4050 4.2520 0.4550 ;
      RECT 4.2310 0.9200 4.6610 0.9700 ;
      RECT 4.6110 0.8310 4.6610 0.9200 ;
      RECT 4.2310 0.9700 4.2810 1.0340 ;
      RECT 4.2310 0.5050 4.2810 0.9200 ;
      RECT 3.9870 1.4200 5.2930 1.4700 ;
      RECT 7.0270 1.1990 8.3250 1.2490 ;
      RECT 7.6350 0.5270 8.2330 0.5770 ;
      RECT 8.1830 0.5770 8.2330 0.7700 ;
      RECT 8.1830 0.3480 8.2330 0.5270 ;
      RECT 7.8790 0.5770 7.9290 0.8870 ;
      RECT 7.8790 0.1260 7.9290 0.5270 ;
      RECT 8.3190 0.1320 8.5530 0.1820 ;
      RECT 7.5750 1.0570 8.0240 1.1070 ;
      RECT 7.5750 0.6770 7.6250 1.0570 ;
      RECT 7.5350 0.6270 7.6250 0.6770 ;
      RECT 7.5350 0.4770 7.5850 0.6270 ;
      RECT 7.5350 0.4270 7.6250 0.4770 ;
      RECT 7.5750 0.1260 7.6250 0.4270 ;
      RECT 2.6190 1.5240 3.7650 1.5740 ;
      RECT 5.6590 0.0880 5.8930 0.1380 ;
      RECT 0.7190 0.5100 1.2570 0.5600 ;
      RECT 1.1750 1.1330 1.5610 1.1830 ;
      RECT 0.7190 0.9410 0.9530 0.9910 ;
      RECT 2.8630 0.7130 2.9890 0.7630 ;
      RECT 2.8630 0.7630 2.9130 1.0330 ;
      RECT 2.9390 0.5630 2.9890 0.7130 ;
      RECT 2.8470 0.5130 2.9890 0.5630 ;
      RECT 4.5190 0.3840 5.1930 0.4340 ;
      RECT 5.1430 0.4340 5.1930 0.5630 ;
      RECT 5.1430 0.2970 5.1930 0.3840 ;
      RECT 4.9910 0.4340 5.0410 0.9670 ;
      RECT 4.9910 0.9670 5.2090 1.0170 ;
      RECT 4.9910 1.0170 5.0410 1.1200 ;
      RECT 4.9910 1.1700 5.0410 1.2700 ;
      RECT 4.5190 1.1200 5.0410 1.1700 ;
      RECT 3.5270 0.9680 4.0390 1.0180 ;
      RECT 3.9860 0.9080 4.0360 0.9680 ;
      RECT 3.9860 0.8580 4.0690 0.9080 ;
      RECT 1.4520 0.6020 1.6370 0.6520 ;
      RECT 0.2050 0.8410 1.5020 0.8910 ;
      RECT 1.4520 0.6520 1.5020 0.8410 ;
      RECT 0.2050 0.5260 0.2550 0.8410 ;
      RECT 0.2790 0.8910 0.3290 1.2140 ;
      RECT 0.2050 0.4760 0.3290 0.5260 ;
      RECT 0.2790 0.3160 0.3290 0.4760 ;
      RECT 5.9630 0.6320 6.5010 0.6820 ;
      RECT 5.2950 0.4500 5.3450 0.5630 ;
      RECT 5.2950 0.2970 5.3450 0.4000 ;
      RECT 5.2960 1.2290 5.3460 1.3530 ;
      RECT 5.6600 0.4500 5.7100 1.1790 ;
      RECT 5.2960 1.1790 5.8170 1.2290 ;
    LAYER PO ;
      RECT 5.5330 0.0660 5.5630 0.6910 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.7090 0.0660 3.7390 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 3.1010 0.8400 3.1310 1.6060 ;
      RECT 5.5330 0.9390 5.5630 1.6060 ;
      RECT 5.2290 0.0660 5.2590 0.6370 ;
      RECT 3.1010 0.0660 3.1310 0.6370 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 4.7730 0.0660 4.8030 0.6910 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 9.3330 0.0660 9.3630 1.6060 ;
      RECT 4.4690 0.8920 4.4990 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 5.2290 0.8390 5.2590 1.6060 ;
      RECT 9.4850 0.0660 9.5150 1.6060 ;
      RECT 9.9410 0.0660 9.9710 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 9.6370 0.0660 9.6670 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 9.7890 0.0660 9.8190 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 3.5570 0.0680 3.5870 0.6180 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 4.4690 0.0660 4.4990 0.6910 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 7.0530 0.0670 7.0830 1.6050 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 4.7730 0.8390 4.8030 1.6060 ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 3.5570 0.7300 3.5870 1.6060 ;
    LAYER NWELL ;
      RECT 7.4080 0.4910 9.4190 1.0830 ;
      RECT -0.1150 1.5430 10.1490 1.7730 ;
      RECT -0.1150 0.6790 6.9460 1.5430 ;
      RECT 9.8790 0.6790 10.1490 1.5430 ;
  END
END RSDFFNSRX2_LVT

MACRO RSDFFNX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.184 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 8.0150 0.9440 9.4820 1.0040 ;
        RECT 9.3720 0.6900 9.4820 0.9440 ;
    END
  END VDDG

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6780 0.7250 0.7280 ;
        RECT 0.4010 0.5510 0.5110 0.6780 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 1.1610 1.0110 1.3160 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 10.1840 0.0300 ;
        RECT 2.2080 0.0300 2.2580 0.3070 ;
        RECT 9.0950 0.0300 9.1450 0.3120 ;
        RECT 8.7910 0.0300 8.8410 0.2020 ;
        RECT 0.5830 0.0300 0.6330 0.5120 ;
        RECT 8.0310 0.0300 8.0810 0.2110 ;
        RECT 1.7990 0.0300 1.8490 0.4050 ;
        RECT 6.9670 0.0300 7.0170 0.2410 ;
        RECT 0.4310 0.0300 0.4810 0.4450 ;
        RECT 1.6470 0.0300 1.6970 0.4210 ;
        RECT 6.7030 0.0300 6.7530 0.2830 ;
        RECT 2.2080 0.3070 3.9770 0.3570 ;
        RECT 4.8230 0.2830 6.7540 0.3330 ;
        RECT 2.2550 0.3570 2.3050 0.5570 ;
        RECT 3.9270 0.3570 3.9770 0.5770 ;
        RECT 3.3190 0.3570 3.3690 0.5580 ;
        RECT 3.4710 0.3570 3.5210 0.5580 ;
        RECT 6.6630 0.3330 6.7130 0.4430 ;
    END
  END VSS

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0740 1.4650 2.2460 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.1190 0.9690 7.6530 1.0190 ;
        RECT 7.1190 1.0190 7.3510 1.1290 ;
        RECT 7.6030 0.3510 7.6530 0.9690 ;
        RECT 7.1190 1.1290 7.1690 1.3270 ;
        RECT 7.1030 0.3010 7.6530 0.3510 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.8150 0.1570 6.8650 0.4010 ;
        RECT 6.8150 0.4010 7.5150 0.4510 ;
        RECT 7.3930 0.4510 7.5150 0.5380 ;
        RECT 7.4650 0.5380 7.5150 0.8590 ;
        RECT 6.8150 0.8590 7.5150 0.9090 ;
        RECT 6.8150 0.9090 6.8650 1.2320 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 10.1840 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 0.4310 1.0130 0.4810 1.6420 ;
        RECT 1.6470 1.1230 1.6970 1.6420 ;
        RECT 1.7990 1.1210 1.8490 1.6420 ;
        RECT 5.0310 1.3400 5.0810 1.6420 ;
        RECT 1.9620 1.3400 2.0120 1.6420 ;
        RECT 1.9620 1.2900 7.0180 1.3400 ;
        RECT 1.9620 1.2670 2.0120 1.2900 ;
        RECT 6.9670 0.9590 7.0170 1.2900 ;
        RECT 4.8390 0.9730 4.8890 1.2900 ;
    END
  END VDD

  PIN RETN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.3370 1.4080 8.7190 1.4580 ;
        RECT 8.6090 1.3130 8.7190 1.4080 ;
    END
    ANTENNAGATEAREA 0.084 ;
  END RETN

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2520 1.3330 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI
  OBS
    LAYER M1 ;
      RECT 1.0230 0.4100 1.3930 0.4600 ;
      RECT 1.0230 1.0200 1.7000 1.0700 ;
      RECT 1.6500 0.7520 1.7000 1.0200 ;
      RECT 1.6500 0.7280 1.7370 0.7520 ;
      RECT 1.6870 0.5520 1.7370 0.6780 ;
      RECT 1.3430 0.5020 1.7370 0.5520 ;
      RECT 9.2470 0.5620 9.5410 0.6120 ;
      RECT 9.3820 0.4120 9.4320 0.5620 ;
      RECT 9.2470 0.3620 9.4320 0.4120 ;
      RECT 9.2470 0.6120 9.2970 0.8340 ;
      RECT 8.0830 0.8340 9.2970 0.8840 ;
      RECT 9.2470 0.1260 9.2970 0.3620 ;
      RECT 8.0830 0.4200 8.1330 0.8340 ;
      RECT 8.0830 0.3700 8.2510 0.4200 ;
      RECT 4.6870 0.5130 4.7770 0.5630 ;
      RECT 4.7270 0.5630 4.7770 0.7670 ;
      RECT 4.6470 0.7670 4.7770 0.8170 ;
      RECT 4.6870 0.3270 4.7370 0.5130 ;
      RECT 4.5350 0.2770 4.7370 0.3270 ;
      RECT 4.6470 0.8170 4.6970 0.9740 ;
      RECT 4.5350 0.3270 4.5850 0.5560 ;
      RECT 4.6470 0.9740 4.7370 1.0240 ;
      RECT 4.6870 1.0240 4.7370 1.1900 ;
      RECT 4.5350 1.1900 4.7370 1.2400 ;
      RECT 4.5350 0.9740 4.5850 1.1900 ;
      RECT 4.9510 0.7670 5.1930 0.8170 ;
      RECT 5.1430 0.8170 5.1930 1.2400 ;
      RECT 4.9510 0.4530 5.0010 0.7670 ;
      RECT 4.8270 0.4030 5.1940 0.4530 ;
      RECT 5.1430 0.4530 5.1930 0.5770 ;
      RECT 4.8270 0.4530 4.8770 0.8670 ;
      RECT 4.7470 0.8670 4.8770 0.9170 ;
      RECT 2.6350 0.6130 2.8530 0.6630 ;
      RECT 2.6350 0.5630 2.6850 0.6130 ;
      RECT 2.6350 0.6630 2.6850 0.7540 ;
      RECT 2.5430 0.5130 2.6850 0.5630 ;
      RECT 2.5420 0.7540 2.6850 0.8040 ;
      RECT 3.7350 0.8670 4.0170 0.9170 ;
      RECT 3.9670 0.9170 4.0170 1.1270 ;
      RECT 3.0150 1.1270 4.0170 1.1770 ;
      RECT 3.0150 1.1770 3.0650 1.2400 ;
      RECT 3.0150 1.0660 3.1150 1.1270 ;
      RECT 3.0650 0.9170 3.1150 1.0660 ;
      RECT 3.0150 0.4130 3.0650 0.8670 ;
      RECT 3.0150 0.8670 3.3090 0.9170 ;
      RECT 3.7350 0.6070 3.7850 0.8670 ;
      RECT 3.7350 0.5570 3.8250 0.6070 ;
      RECT 3.7750 0.4130 3.8250 0.5570 ;
      RECT 0.7190 0.5100 1.2570 0.5600 ;
      RECT 1.9520 0.9670 3.0050 1.0170 ;
      RECT 1.9520 1.0170 2.0020 1.0760 ;
      RECT 1.9520 0.8280 2.0020 0.9670 ;
      RECT 1.9520 0.7780 2.0410 0.8280 ;
      RECT 1.9910 0.6280 2.0410 0.7780 ;
      RECT 1.9520 0.5780 2.0410 0.6280 ;
      RECT 1.9520 0.3190 2.0020 0.5780 ;
      RECT 1.1750 1.1330 1.5610 1.1830 ;
      RECT 0.8870 0.3100 1.5450 0.3600 ;
      RECT 1.4950 0.3600 1.5450 0.3920 ;
      RECT 0.8870 0.3600 0.9370 0.3920 ;
      RECT 8.9430 0.5890 9.1360 0.6390 ;
      RECT 9.0860 0.5120 9.1360 0.5890 ;
      RECT 9.0860 0.4620 9.2370 0.5120 ;
      RECT 9.0860 0.4120 9.1360 0.4620 ;
      RECT 8.9430 0.3620 9.1360 0.4120 ;
      RECT 8.9430 0.6390 8.9930 0.7790 ;
      RECT 8.9430 0.1260 8.9930 0.3620 ;
      RECT 4.4430 0.6130 4.6770 0.6630 ;
      RECT 2.6190 1.5240 4.6770 1.5740 ;
      RECT 2.3150 0.0940 4.3730 0.1440 ;
      RECT 5.3550 0.6130 6.2570 0.6630 ;
      RECT 6.2070 0.3830 6.2570 0.6130 ;
      RECT 5.5590 0.6630 5.6090 0.9670 ;
      RECT 5.5590 0.9670 6.2570 1.0170 ;
      RECT 6.2070 1.0170 6.2570 1.2400 ;
      RECT 8.6390 0.4620 8.9330 0.5120 ;
      RECT 8.6390 0.1820 8.6890 0.4620 ;
      RECT 8.6390 0.5120 8.6890 0.6350 ;
      RECT 8.3190 0.1320 8.6890 0.1820 ;
      RECT 8.3190 0.6350 8.6890 0.6850 ;
      RECT 5.5070 1.5280 9.5430 1.5780 ;
      RECT 5.6590 0.7130 5.8930 0.7630 ;
      RECT 4.2910 0.8670 4.5450 0.9170 ;
      RECT 2.1030 0.6130 2.5490 0.6630 ;
      RECT 2.1030 0.8670 2.8530 0.9170 ;
      RECT 2.1030 0.4130 2.1530 0.6130 ;
      RECT 2.1030 0.6630 2.1530 0.8670 ;
      RECT 0.7190 0.9410 0.9530 0.9910 ;
      RECT 3.8350 0.6670 4.2210 0.7170 ;
      RECT 7.3310 1.2310 8.4770 1.2810 ;
      RECT 6.7910 0.5010 7.0930 0.5510 ;
      RECT 7.0430 0.5510 7.0930 0.6790 ;
      RECT 6.7910 0.5510 6.8410 0.6130 ;
      RECT 6.4190 0.6130 6.8410 0.6630 ;
      RECT 1.4520 0.6020 1.6370 0.6520 ;
      RECT 0.2050 0.8410 1.5020 0.8910 ;
      RECT 1.4520 0.6520 1.5020 0.8410 ;
      RECT 0.2050 0.5260 0.2550 0.8410 ;
      RECT 0.2790 0.8910 0.3290 1.2140 ;
      RECT 0.2050 0.4760 0.3290 0.5260 ;
      RECT 0.2790 0.3160 0.3290 0.4760 ;
      RECT 7.8790 1.0800 8.3250 1.1300 ;
      RECT 7.8790 0.1260 7.9290 1.0800 ;
      RECT 4.4230 0.0920 6.5020 0.1420 ;
      RECT 4.4230 0.1420 4.4730 0.1940 ;
      RECT 4.3830 0.1940 4.4730 0.2440 ;
      RECT 4.3830 0.2440 4.4330 0.5130 ;
      RECT 4.2310 0.5130 4.4330 0.5630 ;
      RECT 4.2310 0.2770 4.2810 0.5130 ;
      RECT 4.2710 0.5630 4.3210 0.7670 ;
      RECT 4.1910 0.7670 4.3210 0.8170 ;
      RECT 4.1910 0.8170 4.2410 0.9670 ;
      RECT 4.1910 0.9670 4.2810 1.0170 ;
      RECT 4.2310 1.0170 4.2810 1.1900 ;
      RECT 4.2310 1.1900 4.4330 1.2400 ;
      RECT 4.3830 0.9740 4.4330 1.1900 ;
      RECT 8.1830 0.4940 8.5370 0.5440 ;
      RECT 8.4870 0.3480 8.5370 0.4940 ;
      RECT 8.1830 0.5440 8.2330 0.7340 ;
      RECT 5.0510 0.6270 5.3050 0.6770 ;
      RECT 5.2550 0.5630 5.3050 0.6270 ;
      RECT 5.2550 0.6770 5.3050 1.0670 ;
      RECT 5.2550 0.5130 6.1210 0.5630 ;
      RECT 5.2550 1.0670 6.1210 1.1170 ;
      RECT 3.3030 0.9670 3.9170 1.0170 ;
      RECT 3.1670 0.4070 3.2170 0.6190 ;
      RECT 3.4710 0.6690 3.5210 0.9670 ;
      RECT 3.1670 0.6190 3.5210 0.6690 ;
      RECT 5.9630 0.7590 7.4130 0.8090 ;
      RECT 6.8910 0.6420 6.9410 0.7590 ;
      RECT 6.5110 0.8090 6.5610 1.2400 ;
      RECT 6.3190 0.5630 6.3690 0.7590 ;
      RECT 6.3190 0.5130 6.5610 0.5630 ;
      RECT 6.5110 0.3830 6.5610 0.5130 ;
      RECT 1.6500 0.7020 1.9410 0.7280 ;
      RECT 1.6870 0.6780 1.9410 0.7020 ;
      RECT 1.3430 0.4600 1.3930 0.5020 ;
    LAYER PO ;
      RECT 9.7890 0.0660 9.8190 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 9.4850 0.0660 9.5150 1.6060 ;
      RECT 5.8370 0.0660 5.8670 0.7910 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 9.6370 0.0660 9.6670 1.6060 ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 4.4690 0.0660 4.4990 0.6910 ;
      RECT 4.0130 0.0660 4.0430 0.6370 ;
      RECT 2.7970 0.8390 2.8270 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 5.8370 0.9390 5.8670 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 3.7090 0.0660 3.7390 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 4.4690 0.8390 4.4990 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 9.3330 0.0660 9.3630 1.6060 ;
      RECT 5.3810 0.9590 5.4110 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 7.3570 0.0670 7.3870 1.6050 ;
      RECT 3.5570 0.9390 3.5870 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 3.5570 0.0660 3.5870 0.6370 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 2.7970 0.0660 2.8270 0.6910 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 10.0930 0.0660 10.1230 1.6060 ;
      RECT 4.0130 0.9390 4.0430 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 9.9410 0.0660 9.9710 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 5.3810 0.0660 5.4110 0.6910 ;
    LAYER NWELL ;
      RECT -0.1160 1.5430 10.2940 1.7730 ;
      RECT -0.1160 0.6790 7.2510 1.5430 ;
      RECT 10.0190 0.6790 10.2940 1.5430 ;
      RECT 7.7130 0.4910 9.5590 1.0830 ;
  END
END RSDFFNX1_LVT

MACRO RSDFFNX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.488 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.2710 0.2710 7.9690 0.3210 ;
        RECT 7.8510 0.3210 7.9690 0.3590 ;
        RECT 7.8510 0.2500 7.9690 0.2710 ;
        RECT 7.2710 0.1490 7.3210 0.2710 ;
        RECT 7.9190 0.3590 7.9690 0.9330 ;
        RECT 7.8510 0.2490 7.9610 0.2500 ;
        RECT 7.2710 0.9330 7.9690 0.9830 ;
        RECT 7.2710 0.9830 7.3210 1.2240 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 8.3190 0.9540 9.7860 1.0140 ;
        RECT 9.6760 0.6900 9.7860 0.9540 ;
    END
  END VDDG

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.9670 0.1490 7.0170 0.4020 ;
        RECT 6.9670 0.4020 7.8190 0.4520 ;
        RECT 7.6970 0.4520 7.8190 0.5120 ;
        RECT 7.7690 0.5120 7.8190 0.8330 ;
        RECT 6.9670 0.8330 7.8190 0.8830 ;
        RECT 6.9670 0.8830 7.0170 1.2240 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6780 0.7250 0.7280 ;
        RECT 0.4010 0.5510 0.5110 0.6780 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 1.1610 1.0110 1.3160 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 10.4880 0.0300 ;
        RECT 2.2080 0.0300 2.2580 0.3070 ;
        RECT 9.3990 0.0300 9.4490 0.3120 ;
        RECT 0.4310 0.0300 0.4810 0.4340 ;
        RECT 1.6470 0.0300 1.6970 0.4050 ;
        RECT 9.0950 0.0300 9.1450 0.2020 ;
        RECT 0.5830 0.0300 0.6330 0.5120 ;
        RECT 7.4230 0.0300 7.4730 0.2210 ;
        RECT 8.3350 0.0300 8.3850 0.2060 ;
        RECT 6.8150 0.0300 6.8650 0.4090 ;
        RECT 1.7990 0.0300 1.8490 0.4050 ;
        RECT 7.1190 0.0300 7.1690 0.3200 ;
        RECT 6.7030 0.0300 6.7530 0.2830 ;
        RECT 2.2080 0.3070 3.9770 0.3570 ;
        RECT 4.8230 0.2830 6.7540 0.3330 ;
        RECT 2.2550 0.3570 2.3050 0.5570 ;
        RECT 3.9270 0.3570 3.9770 0.5770 ;
        RECT 3.3190 0.3570 3.3690 0.5580 ;
        RECT 3.4710 0.3570 3.5210 0.5580 ;
        RECT 6.6630 0.3330 6.7130 0.4430 ;
    END
  END VSS

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0740 1.4650 2.2460 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 10.4880 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 1.7990 1.1310 1.8490 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 1.6470 1.1310 1.6970 1.6420 ;
        RECT 5.0310 1.3400 5.0810 1.6420 ;
        RECT 1.9620 1.3400 2.0120 1.6420 ;
        RECT 1.9620 1.2900 7.4730 1.3400 ;
        RECT 7.4230 1.0530 7.4730 1.2900 ;
        RECT 7.1190 0.9610 7.1690 1.2900 ;
        RECT 6.8150 0.9130 6.8650 1.2900 ;
        RECT 4.8390 0.9730 4.8890 1.2900 ;
    END
  END VDD

  PIN RETN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.3370 1.4080 9.0230 1.4580 ;
        RECT 8.9130 1.3130 9.0230 1.4080 ;
    END
    ANTENNAGATEAREA 0.084 ;
  END RETN

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2520 1.3330 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI
  OBS
    LAYER M1 ;
      RECT 5.9630 0.7130 7.7170 0.7630 ;
      RECT 6.5110 0.7630 6.5610 1.2400 ;
      RECT 6.3190 0.5630 6.3690 0.7130 ;
      RECT 6.3190 0.5130 6.5610 0.5630 ;
      RECT 6.5110 0.3830 6.5610 0.5130 ;
      RECT 6.8910 0.6420 6.9410 0.7130 ;
      RECT 7.0430 0.6420 7.0930 0.7130 ;
      RECT 5.5070 1.5280 9.8470 1.5780 ;
      RECT 5.6590 0.7130 5.8930 0.7630 ;
      RECT 9.3900 0.4120 9.4400 0.4620 ;
      RECT 9.3900 0.4620 9.5410 0.5120 ;
      RECT 9.3900 0.5120 9.4400 0.5890 ;
      RECT 9.2470 0.5890 9.4400 0.6390 ;
      RECT 9.2470 0.3620 9.4400 0.4120 ;
      RECT 9.2470 0.1260 9.2970 0.3620 ;
      RECT 9.2470 0.6390 9.2970 0.7650 ;
      RECT 4.6870 0.5130 4.7770 0.5630 ;
      RECT 4.7270 0.5630 4.7770 0.7670 ;
      RECT 4.6470 0.7670 4.7770 0.8170 ;
      RECT 4.5350 0.3270 4.5850 0.5560 ;
      RECT 4.5350 0.2770 4.7370 0.3270 ;
      RECT 4.6870 0.3270 4.7370 0.5130 ;
      RECT 4.6470 0.8170 4.6970 0.9740 ;
      RECT 4.6470 0.9740 4.7370 1.0240 ;
      RECT 4.6870 1.0240 4.7370 1.1900 ;
      RECT 4.5350 1.1900 4.7370 1.2400 ;
      RECT 4.5350 0.9740 4.5850 1.1900 ;
      RECT 5.0510 0.6270 5.3050 0.6770 ;
      RECT 5.2550 0.5630 5.3050 0.6270 ;
      RECT 5.2550 0.6770 5.3050 1.0670 ;
      RECT 5.2550 0.5130 6.1210 0.5630 ;
      RECT 5.2550 1.0670 6.1210 1.1170 ;
      RECT 3.3030 0.9670 3.9170 1.0170 ;
      RECT 3.1670 0.4070 3.2170 0.6190 ;
      RECT 3.4710 0.6690 3.5210 0.9670 ;
      RECT 3.1670 0.6190 3.5210 0.6690 ;
      RECT 1.6500 0.7020 1.9410 0.7280 ;
      RECT 1.6870 0.6780 1.9410 0.7020 ;
      RECT 1.3430 0.4600 1.3930 0.5020 ;
      RECT 1.0230 0.4100 1.3930 0.4600 ;
      RECT 1.0230 1.0200 1.7000 1.0700 ;
      RECT 1.6500 0.7520 1.7000 1.0200 ;
      RECT 1.6500 0.7280 1.7370 0.7520 ;
      RECT 1.6870 0.5520 1.7370 0.6780 ;
      RECT 1.3430 0.5020 1.7370 0.5520 ;
      RECT 9.5510 0.5620 9.8450 0.6120 ;
      RECT 9.6860 0.4120 9.7360 0.5620 ;
      RECT 9.5510 0.3620 9.7360 0.4120 ;
      RECT 9.5510 0.6120 9.6010 0.8330 ;
      RECT 8.3870 0.8330 9.6010 0.8830 ;
      RECT 9.5510 0.1260 9.6010 0.3620 ;
      RECT 8.3870 0.4200 8.4370 0.8330 ;
      RECT 8.3870 0.3700 8.5550 0.4200 ;
      RECT 4.9510 0.7670 5.1930 0.8170 ;
      RECT 5.1430 0.8170 5.1930 1.2400 ;
      RECT 4.9510 0.4530 5.0010 0.7670 ;
      RECT 4.8270 0.4030 5.1940 0.4530 ;
      RECT 5.1430 0.4530 5.1930 0.5770 ;
      RECT 4.8270 0.4530 4.8770 0.8670 ;
      RECT 4.7470 0.8670 4.8770 0.9170 ;
      RECT 2.1030 0.6130 2.5490 0.6630 ;
      RECT 2.1030 0.8670 2.8530 0.9170 ;
      RECT 2.1030 0.4130 2.1530 0.6130 ;
      RECT 2.1030 0.6630 2.1530 0.8670 ;
      RECT 0.8870 0.3100 1.5450 0.3600 ;
      RECT 0.8870 0.3600 0.9370 0.3920 ;
      RECT 1.4950 0.3600 1.5450 0.3920 ;
      RECT 7.6350 1.2000 8.7810 1.2500 ;
      RECT 5.3550 0.6130 6.2570 0.6630 ;
      RECT 6.2070 0.3830 6.2570 0.6130 ;
      RECT 5.5590 0.6630 5.6090 0.9670 ;
      RECT 5.5590 0.9670 6.2570 1.0170 ;
      RECT 6.2070 1.0170 6.2570 1.2400 ;
      RECT 2.6350 0.6130 2.8530 0.6630 ;
      RECT 2.6350 0.5630 2.6850 0.6130 ;
      RECT 2.6350 0.6630 2.6850 0.7540 ;
      RECT 2.5430 0.5130 2.6850 0.5630 ;
      RECT 2.5420 0.7540 2.6850 0.8040 ;
      RECT 3.7350 0.8670 4.0170 0.9170 ;
      RECT 3.9670 0.9170 4.0170 1.1270 ;
      RECT 3.0150 1.1270 4.0170 1.1770 ;
      RECT 3.0150 1.1770 3.0650 1.2400 ;
      RECT 3.0150 1.0660 3.1150 1.1270 ;
      RECT 3.0650 0.9170 3.1150 1.0660 ;
      RECT 3.0150 0.4130 3.0650 0.8670 ;
      RECT 3.0150 0.8670 3.3090 0.9170 ;
      RECT 3.7350 0.6070 3.7850 0.8670 ;
      RECT 3.7350 0.5570 3.8250 0.6070 ;
      RECT 3.7750 0.4130 3.8250 0.5570 ;
      RECT 0.7190 0.5100 1.2570 0.5600 ;
      RECT 1.9520 0.9670 3.0050 1.0170 ;
      RECT 1.9520 1.0170 2.0020 1.0760 ;
      RECT 1.9520 0.8280 2.0020 0.9670 ;
      RECT 1.9520 0.7780 2.0410 0.8280 ;
      RECT 1.9910 0.6280 2.0410 0.7780 ;
      RECT 1.9520 0.5780 2.0410 0.6280 ;
      RECT 1.9520 0.3190 2.0020 0.5780 ;
      RECT 1.1750 1.1330 1.5610 1.1830 ;
      RECT 4.4430 0.6130 4.6770 0.6630 ;
      RECT 2.6190 1.5240 4.6770 1.5740 ;
      RECT 2.3150 0.0940 4.3730 0.1440 ;
      RECT 4.2910 0.8670 4.5450 0.9170 ;
      RECT 0.7190 0.9410 0.9530 0.9910 ;
      RECT 3.8350 0.6670 4.2210 0.7170 ;
      RECT 6.4190 0.6130 6.7870 0.6630 ;
      RECT 6.7370 0.5700 6.7870 0.6130 ;
      RECT 6.7370 0.5200 7.2270 0.5700 ;
      RECT 7.1770 0.5700 7.2270 0.6040 ;
      RECT 7.1770 0.6040 7.4130 0.6540 ;
      RECT 1.4520 0.6020 1.6370 0.6520 ;
      RECT 0.2050 0.8410 1.5020 0.8910 ;
      RECT 1.4520 0.6520 1.5020 0.8410 ;
      RECT 0.2050 0.5260 0.2550 0.8410 ;
      RECT 0.2790 0.8910 0.3290 1.2140 ;
      RECT 0.2050 0.4760 0.3290 0.5260 ;
      RECT 0.2790 0.3160 0.3290 0.4760 ;
      RECT 8.1830 1.0860 8.6290 1.1360 ;
      RECT 8.1830 0.1260 8.2330 1.0860 ;
      RECT 4.4230 0.0920 6.5020 0.1420 ;
      RECT 4.4230 0.1420 4.4730 0.1940 ;
      RECT 4.3830 0.1940 4.4730 0.2440 ;
      RECT 4.3830 0.2440 4.4330 0.5130 ;
      RECT 4.2310 0.5130 4.4330 0.5630 ;
      RECT 4.2310 0.2770 4.2810 0.5130 ;
      RECT 4.2710 0.5630 4.3210 0.7670 ;
      RECT 4.1910 0.7670 4.3210 0.8170 ;
      RECT 4.1910 0.8170 4.2410 0.9670 ;
      RECT 4.1910 0.9670 4.2810 1.0170 ;
      RECT 4.2310 1.0170 4.2810 1.1900 ;
      RECT 4.2310 1.1900 4.4330 1.2400 ;
      RECT 4.3830 0.9740 4.4330 1.1900 ;
      RECT 8.4870 0.4940 8.8410 0.5440 ;
      RECT 8.7910 0.3480 8.8410 0.4940 ;
      RECT 8.4870 0.5440 8.5370 0.7600 ;
      RECT 8.9430 0.4620 9.2370 0.5120 ;
      RECT 8.9430 0.5120 8.9930 0.6350 ;
      RECT 8.9430 0.1820 8.9930 0.4620 ;
      RECT 8.6230 0.6350 8.9930 0.6850 ;
      RECT 8.6230 0.1320 8.9930 0.1820 ;
    LAYER PO ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 10.3970 0.0660 10.4270 1.6060 ;
      RECT 4.0130 0.9390 4.0430 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 10.2450 0.0660 10.2750 1.6060 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 5.3810 0.0660 5.4110 0.6910 ;
      RECT 10.0930 0.0660 10.1230 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 9.7890 0.0660 9.8190 1.6060 ;
      RECT 5.8370 0.0660 5.8670 0.7910 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 9.9410 0.0660 9.9710 1.6060 ;
      RECT 9.4850 0.0660 9.5150 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 4.4690 0.0660 4.4990 0.6910 ;
      RECT 4.0130 0.0660 4.0430 0.6370 ;
      RECT 2.7970 0.8390 2.8270 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 5.8370 0.9390 5.8670 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 3.7090 0.0660 3.7390 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 4.4690 0.8390 4.4990 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 9.3330 0.0660 9.3630 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 9.6370 0.0660 9.6670 1.6060 ;
      RECT 5.3810 0.9590 5.4110 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 7.6610 0.0670 7.6910 1.6050 ;
      RECT 3.5570 0.9390 3.5870 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 3.5570 0.0660 3.5870 0.6370 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 2.7970 0.0660 2.8270 0.6910 ;
    LAYER NWELL ;
      RECT -0.1160 1.5430 10.5980 1.7730 ;
      RECT -0.1160 0.6790 7.5550 1.5430 ;
      RECT 10.3230 0.6790 10.5980 1.5430 ;
      RECT 8.0170 0.4910 9.8630 1.0830 ;
  END
END RSDFFNX2_LVT

MACRO RSDFFSRARX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.032 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 10.0320 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 2.1030 1.1310 2.1530 1.6420 ;
        RECT 1.7990 1.1310 1.8490 1.6420 ;
        RECT 1.6470 1.1310 1.6970 1.6420 ;
        RECT 2.7110 1.2940 2.7610 1.6420 ;
        RECT 3.9670 1.2700 4.0170 1.6420 ;
        RECT 8.0710 1.4540 8.1210 1.6420 ;
        RECT 2.5390 1.2440 2.7610 1.2940 ;
        RECT 3.7580 1.2200 4.9050 1.2700 ;
        RECT 5.5990 1.4040 8.1210 1.4540 ;
        RECT 5.5990 1.2790 5.6490 1.4040 ;
        RECT 6.6630 0.9590 6.7130 1.4040 ;
        RECT 6.2070 0.9530 6.2570 1.4040 ;
    END
  END VDD

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.5110 0.4010 7.2110 0.4510 ;
        RECT 6.5110 0.1570 6.5610 0.4010 ;
        RECT 7.0890 0.4510 7.2110 0.5380 ;
        RECT 7.1610 0.5380 7.2110 0.8590 ;
        RECT 6.5110 0.8590 7.2110 0.9090 ;
        RECT 6.5110 0.9090 6.5610 1.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.8150 0.9690 7.3490 1.0190 ;
        RECT 7.2990 0.3510 7.3490 0.9690 ;
        RECT 6.8150 1.0190 7.0470 1.1290 ;
        RECT 6.7990 0.3010 7.3490 0.3510 ;
        RECT 6.8150 1.1290 6.8650 1.3270 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4670 1.4650 2.6390 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 10.0320 0.0300 ;
        RECT 2.1030 0.0300 2.1530 0.2970 ;
        RECT 9.0950 0.0300 9.1450 0.4260 ;
        RECT 1.6470 0.0300 1.6970 0.4050 ;
        RECT 6.6630 0.0300 6.7130 0.2410 ;
        RECT 1.7990 0.0300 1.8490 0.4050 ;
        RECT 7.7270 0.0300 7.7770 0.4260 ;
        RECT 0.5830 0.0300 0.6330 0.5120 ;
        RECT 0.4310 0.0300 0.4810 0.4340 ;
        RECT 8.6390 0.0300 8.6890 0.1980 ;
        RECT 6.3830 0.0300 6.4330 0.3000 ;
        RECT 2.1030 0.2970 3.9770 0.3470 ;
        RECT 5.5830 0.3000 6.4330 0.3500 ;
        RECT 3.7750 0.3470 3.8250 0.5570 ;
        RECT 2.5590 0.3470 2.6090 0.5570 ;
        RECT 2.7110 0.3470 2.7610 0.5570 ;
        RECT 2.1030 0.3470 2.1530 0.4050 ;
        RECT 3.9270 0.2380 3.9770 0.2970 ;
        RECT 3.9270 0.1880 4.9050 0.2380 ;
        RECT 4.2310 0.2380 4.2810 0.3490 ;
    END
  END VSS

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4390 0.0970 5.6890 0.1380 ;
        RECT 3.4390 0.1380 3.5970 0.2100 ;
        RECT 5.6390 0.1380 5.6890 0.2000 ;
        RECT 3.5470 0.0880 5.6890 0.0970 ;
        RECT 5.6390 0.2000 6.1810 0.2500 ;
        RECT 6.1310 0.0880 6.1810 0.2000 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.2170 0.2490 9.3270 0.3590 ;
        RECT 9.2280 0.3590 9.2780 0.5270 ;
        RECT 9.0030 0.5270 9.2780 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.5050 0.7050 4.6610 0.7310 ;
        RECT 4.5050 0.7310 4.9650 0.7810 ;
        RECT 4.6110 0.5970 4.6610 0.7050 ;
        RECT 4.5050 0.7810 4.6610 0.8150 ;
        RECT 4.9150 0.7810 4.9650 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 7.7110 0.9480 9.3290 1.0080 ;
        RECT 9.2190 0.6900 9.3290 0.9480 ;
        RECT 9.0950 0.6270 9.1450 0.9480 ;
    END
  END VDDG

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2520 1.3330 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6780 0.7250 0.7280 ;
        RECT 0.4010 0.5510 0.5110 0.6780 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 1.1610 1.0110 1.3160 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D
  OBS
    LAYER M1 ;
      RECT 5.1430 1.1700 5.1930 1.2700 ;
      RECT 4.6710 1.1200 5.1930 1.1700 ;
      RECT 4.1210 0.8580 4.2210 0.9080 ;
      RECT 4.1210 0.9080 4.1710 0.9680 ;
      RECT 3.6830 0.9680 4.1710 1.0180 ;
      RECT 1.4520 0.6020 1.6370 0.6520 ;
      RECT 0.2050 0.8410 1.5020 0.8910 ;
      RECT 1.4520 0.6520 1.5020 0.8410 ;
      RECT 0.2050 0.5260 0.2550 0.8410 ;
      RECT 0.2790 0.8910 0.3290 1.2140 ;
      RECT 0.2050 0.4760 0.3290 0.5260 ;
      RECT 0.2790 0.3160 0.3290 0.4760 ;
      RECT 3.1670 0.8540 4.0690 0.9040 ;
      RECT 3.1670 0.6130 3.2170 0.8540 ;
      RECT 3.1670 0.9040 3.2170 1.0590 ;
      RECT 3.1670 0.5630 3.3690 0.6130 ;
      RECT 3.1670 1.0590 3.5370 1.1090 ;
      RECT 3.3190 0.4070 3.3690 0.5630 ;
      RECT 3.1670 0.4130 3.2170 0.5630 ;
      RECT 3.1670 1.1090 3.2170 1.3370 ;
      RECT 6.2830 0.6420 6.6370 0.6920 ;
      RECT 6.5870 0.5970 6.6370 0.6420 ;
      RECT 5.8180 0.7290 6.0050 0.7790 ;
      RECT 5.9550 0.7790 6.0050 1.1790 ;
      RECT 5.8180 0.4500 5.8680 0.7290 ;
      RECT 5.4480 1.1790 6.0050 1.2290 ;
      RECT 6.2830 0.4500 6.3330 0.6420 ;
      RECT 5.4470 0.4000 6.3330 0.4500 ;
      RECT 5.4480 1.2290 5.4980 1.3530 ;
      RECT 5.4470 0.4500 5.4970 0.5630 ;
      RECT 5.4470 0.2970 5.4970 0.4000 ;
      RECT 2.9990 0.4120 3.1050 0.4620 ;
      RECT 3.0550 0.4620 3.1050 0.8130 ;
      RECT 3.0150 0.8130 3.1050 0.8630 ;
      RECT 3.0150 0.8630 3.0650 1.0830 ;
      RECT 2.2550 1.0830 3.0650 1.1330 ;
      RECT 3.0150 1.1330 3.0650 1.3540 ;
      RECT 2.2550 0.7520 2.3050 1.0830 ;
      RECT 2.2550 0.7020 2.3450 0.7520 ;
      RECT 2.2950 0.5510 2.3450 0.7020 ;
      RECT 2.2550 0.5010 2.3450 0.5510 ;
      RECT 2.2550 0.4070 2.3050 0.5010 ;
      RECT 2.4070 0.6130 2.8530 0.6630 ;
      RECT 2.4070 0.6630 2.4570 1.0040 ;
      RECT 2.4070 0.4130 2.4570 0.6130 ;
      RECT 2.6180 0.0940 3.3150 0.1440 ;
      RECT 8.0150 0.8200 8.5630 0.8700 ;
      RECT 1.6500 0.7020 1.9410 0.7280 ;
      RECT 1.6870 0.6780 1.9410 0.7020 ;
      RECT 1.3430 0.4600 1.3930 0.5020 ;
      RECT 1.0230 0.4100 1.3930 0.4600 ;
      RECT 1.0230 1.0200 1.7000 1.0700 ;
      RECT 1.6500 0.7520 1.7000 1.0200 ;
      RECT 1.6500 0.7280 1.7370 0.7520 ;
      RECT 1.6870 0.5520 1.7370 0.6780 ;
      RECT 1.3430 0.5020 1.7370 0.5520 ;
      RECT 0.8870 0.3100 1.5450 0.3600 ;
      RECT 1.4950 0.3600 1.5450 0.3920 ;
      RECT 0.8870 0.3600 0.9370 0.3920 ;
      RECT 5.5070 0.8660 5.6560 0.9160 ;
      RECT 5.6060 0.9160 5.6560 0.9670 ;
      RECT 5.6060 0.9670 5.7410 1.0170 ;
      RECT 6.6870 0.6130 7.1090 0.6630 ;
      RECT 6.0550 0.8090 6.1050 1.3010 ;
      RECT 6.0550 0.6780 6.1050 0.7590 ;
      RECT 5.9630 0.6280 6.1050 0.6780 ;
      RECT 6.0550 0.5000 6.1050 0.6280 ;
      RECT 6.3590 0.8090 6.4090 1.3010 ;
      RECT 6.6870 0.6630 6.7370 0.7590 ;
      RECT 6.0550 0.7590 6.7370 0.8090 ;
      RECT 1.9910 0.6280 2.2450 0.6520 ;
      RECT 1.9520 0.6020 2.2450 0.6280 ;
      RECT 1.9910 0.6520 2.0410 0.7780 ;
      RECT 1.9520 0.5780 2.0410 0.6020 ;
      RECT 1.9520 0.7780 2.0410 0.8280 ;
      RECT 1.9520 0.3190 2.0020 0.5780 ;
      RECT 1.9520 0.8280 2.0020 1.0760 ;
      RECT 8.3190 0.7090 8.8570 0.7590 ;
      RECT 4.5190 0.4880 5.0810 0.5380 ;
      RECT 5.0310 0.5380 5.0810 1.0200 ;
      RECT 4.5350 1.0200 5.0810 1.0700 ;
      RECT 4.2710 0.7880 4.3210 1.1200 ;
      RECT 3.3740 0.7380 4.3230 0.7880 ;
      RECT 4.0790 0.5050 4.1290 0.7380 ;
      RECT 4.5350 1.0700 4.5850 1.1200 ;
      RECT 4.0580 1.1200 4.5850 1.1700 ;
      RECT 8.9430 0.6770 8.9930 0.7680 ;
      RECT 8.9030 0.4270 8.9930 0.4620 ;
      RECT 8.9430 0.1260 8.9930 0.4270 ;
      RECT 8.9030 0.6270 8.9930 0.6770 ;
      RECT 8.9030 0.5120 8.9530 0.6270 ;
      RECT 8.6990 0.4770 8.9530 0.5120 ;
      RECT 8.6990 0.4620 8.9930 0.4770 ;
      RECT 4.2910 1.5200 4.9810 1.5700 ;
      RECT 4.7460 0.6130 4.9810 0.6630 ;
      RECT 5.2950 0.8670 5.4370 0.9170 ;
      RECT 5.2950 0.6630 5.3450 0.8670 ;
      RECT 5.2950 0.6130 5.7410 0.6630 ;
      RECT 4.3830 0.9200 4.8130 0.9700 ;
      RECT 4.7630 0.8310 4.8130 0.9200 ;
      RECT 4.3830 0.9700 4.4330 1.0340 ;
      RECT 4.3830 0.5050 4.4330 0.9200 ;
      RECT 4.1390 1.4200 5.4450 1.4700 ;
      RECT 3.3030 1.1900 3.6890 1.2400 ;
      RECT 3.2270 1.3890 3.7650 1.4390 ;
      RECT 4.9950 0.1880 5.5890 0.2380 ;
      RECT 4.9950 0.2380 5.0450 0.2880 ;
      RECT 4.3540 0.2880 5.0450 0.3380 ;
      RECT 3.9470 0.4550 3.9970 0.6130 ;
      RECT 3.6830 0.6130 3.9970 0.6630 ;
      RECT 4.3540 0.3380 4.4040 0.4050 ;
      RECT 3.9470 0.4050 4.4040 0.4550 ;
      RECT 7.0270 1.2120 8.3250 1.2620 ;
      RECT 8.3190 0.1320 8.5530 0.1820 ;
      RECT 7.5750 1.0700 8.0240 1.1200 ;
      RECT 7.5750 0.6770 7.6250 1.0700 ;
      RECT 7.5350 0.6270 7.6250 0.6770 ;
      RECT 7.5350 0.4770 7.5850 0.6270 ;
      RECT 7.5350 0.4270 7.6250 0.4770 ;
      RECT 7.5750 0.1260 7.6250 0.4270 ;
      RECT 2.9230 1.5240 3.9170 1.5740 ;
      RECT 7.6350 0.5270 8.2330 0.5770 ;
      RECT 7.8790 0.5770 7.9290 0.8870 ;
      RECT 7.8790 0.1260 7.9290 0.5270 ;
      RECT 8.1830 0.5770 8.2330 0.7700 ;
      RECT 8.1830 0.3480 8.2330 0.5270 ;
      RECT 5.8110 0.0940 6.0450 0.1440 ;
      RECT 0.7190 0.5100 1.2570 0.5600 ;
      RECT 1.1750 1.1330 1.5610 1.1830 ;
      RECT 0.7190 0.9410 0.9530 0.9910 ;
      RECT 8.5470 1.0870 9.0850 1.1370 ;
      RECT 8.0150 0.2480 8.8570 0.2980 ;
      RECT 5.0490 1.5200 8.0210 1.5700 ;
      RECT 2.8630 0.7130 2.9890 0.7630 ;
      RECT 2.8630 0.7630 2.9130 1.0330 ;
      RECT 2.9390 0.5630 2.9890 0.7130 ;
      RECT 2.8470 0.5130 2.9890 0.5630 ;
      RECT 4.6710 0.3880 5.3450 0.4380 ;
      RECT 5.2950 0.4380 5.3450 0.5630 ;
      RECT 5.2950 0.2970 5.3450 0.3880 ;
      RECT 5.1430 0.4380 5.1930 0.9670 ;
      RECT 5.1430 0.9670 5.3610 1.0170 ;
      RECT 5.1430 1.0170 5.1930 1.1200 ;
    LAYER PO ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 5.6850 0.0660 5.7150 0.6910 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 3.1010 0.8400 3.1310 1.6060 ;
      RECT 5.6850 0.9390 5.7150 1.6060 ;
      RECT 5.3810 0.0660 5.4110 0.6370 ;
      RECT 3.1010 0.0660 3.1310 0.6370 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 3.7090 0.0660 3.7390 0.6910 ;
      RECT 4.9250 0.0660 4.9550 0.6910 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 9.3330 0.0660 9.3630 1.6060 ;
      RECT 4.6210 0.8920 4.6510 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 5.3810 0.8390 5.4110 1.6060 ;
      RECT 9.4850 0.0660 9.5150 1.6060 ;
      RECT 9.9410 0.0660 9.9710 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 9.6370 0.0660 9.6670 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 9.7890 0.0660 9.8190 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 4.6210 0.0660 4.6510 0.6910 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 3.7090 0.9390 3.7390 1.6060 ;
      RECT 7.0530 0.0670 7.0830 1.6050 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 4.9250 0.8390 4.9550 1.6060 ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
    LAYER NWELL ;
      RECT 7.4080 0.4910 9.4190 1.0830 ;
      RECT -0.1150 1.5430 10.1540 1.7730 ;
      RECT -0.1150 0.6790 6.9460 1.5430 ;
      RECT 9.8790 0.6790 10.1540 1.5430 ;
  END
END RSDFFSRARX1_LVT

MACRO RSDFFSRARX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.336 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 10.3360 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 2.1030 1.1310 2.1530 1.6420 ;
        RECT 1.7990 1.1310 1.8490 1.6420 ;
        RECT 1.6470 1.1310 1.6970 1.6420 ;
        RECT 8.3750 1.4540 8.4250 1.6420 ;
        RECT 2.7110 1.2940 2.7610 1.6420 ;
        RECT 3.9670 1.2700 4.0170 1.6420 ;
        RECT 5.5990 1.4040 8.4250 1.4540 ;
        RECT 2.5390 1.2440 2.7610 1.2940 ;
        RECT 3.7580 1.2200 4.9050 1.2700 ;
        RECT 5.5990 1.2790 5.6490 1.4040 ;
        RECT 6.2070 0.9530 6.2570 1.4040 ;
        RECT 7.1190 1.0530 7.1690 1.4040 ;
        RECT 6.5110 0.9130 6.5610 1.4040 ;
        RECT 6.8150 0.9610 6.8650 1.4040 ;
    END
  END VDD

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4670 1.4650 2.6390 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 10.3360 0.0300 ;
        RECT 2.1030 0.0300 2.1530 0.2970 ;
        RECT 6.5110 0.0300 6.5610 0.4090 ;
        RECT 6.8150 0.0300 6.8650 0.3200 ;
        RECT 7.1190 0.0300 7.1690 0.2210 ;
        RECT 9.3990 0.0300 9.4490 0.4260 ;
        RECT 1.6470 0.0300 1.6970 0.4050 ;
        RECT 1.7990 0.0300 1.8490 0.4050 ;
        RECT 8.0310 0.0300 8.0810 0.4260 ;
        RECT 0.5830 0.0300 0.6330 0.5120 ;
        RECT 0.4310 0.0300 0.4810 0.4340 ;
        RECT 8.9430 0.0300 8.9930 0.1980 ;
        RECT 6.3830 0.0300 6.4330 0.3000 ;
        RECT 2.1030 0.2970 3.9770 0.3470 ;
        RECT 5.5830 0.3000 6.4330 0.3500 ;
        RECT 3.7750 0.3470 3.8250 0.5570 ;
        RECT 2.5590 0.3470 2.6090 0.5570 ;
        RECT 2.7110 0.3470 2.7610 0.5570 ;
        RECT 2.1030 0.3470 2.1530 0.4050 ;
        RECT 3.9270 0.2380 3.9770 0.2970 ;
        RECT 3.9270 0.1880 4.9050 0.2380 ;
        RECT 4.2310 0.2380 4.2810 0.3490 ;
    END
  END VSS

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4390 0.0970 5.6890 0.1380 ;
        RECT 3.4390 0.1380 3.5970 0.2100 ;
        RECT 5.6390 0.1380 5.6890 0.2000 ;
        RECT 3.5470 0.0880 5.6890 0.0970 ;
        RECT 5.6390 0.2000 6.1810 0.2500 ;
        RECT 6.1310 0.0880 6.1810 0.2000 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.6630 0.1490 6.7130 0.4020 ;
        RECT 6.6630 0.4020 7.5150 0.4520 ;
        RECT 7.3930 0.4520 7.5150 0.5120 ;
        RECT 7.4650 0.5120 7.5150 0.8430 ;
        RECT 6.6630 0.8430 7.5150 0.8930 ;
        RECT 6.6630 0.8930 6.7130 1.3190 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.5210 0.2490 9.6310 0.3590 ;
        RECT 9.5320 0.3590 9.5820 0.5270 ;
        RECT 9.3070 0.5270 9.5820 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.5050 0.7050 4.6610 0.7310 ;
        RECT 4.5050 0.7310 4.9650 0.7810 ;
        RECT 4.6110 0.5970 4.6610 0.7050 ;
        RECT 4.5050 0.7810 4.6610 0.8150 ;
        RECT 4.9150 0.7810 4.9650 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.5470 0.3210 7.6650 0.3590 ;
        RECT 6.9670 0.2710 7.6650 0.3210 ;
        RECT 7.6150 0.3590 7.6650 0.9430 ;
        RECT 7.5470 0.2490 7.6650 0.2710 ;
        RECT 6.9670 0.1490 7.0170 0.2710 ;
        RECT 6.9670 0.9430 7.6650 0.9930 ;
        RECT 6.9670 0.9930 7.0170 1.3270 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 8.0150 0.9500 9.6330 1.0100 ;
        RECT 9.5230 0.6900 9.6330 0.9500 ;
        RECT 9.3990 0.6270 9.4490 0.9500 ;
    END
  END VDDG

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2520 1.3330 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6780 0.7250 0.7280 ;
        RECT 0.4010 0.5510 0.5110 0.6780 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 1.1610 1.0110 1.3160 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D
  OBS
    LAYER M1 ;
      RECT 5.1430 1.0170 5.1930 1.1200 ;
      RECT 5.1430 1.1700 5.1930 1.2700 ;
      RECT 4.6710 1.1200 5.1930 1.1700 ;
      RECT 4.1210 0.8580 4.2210 0.9080 ;
      RECT 4.1210 0.9080 4.1710 0.9680 ;
      RECT 3.6830 0.9680 4.1710 1.0180 ;
      RECT 1.4520 0.6020 1.6370 0.6520 ;
      RECT 0.2050 0.8410 1.5020 0.8910 ;
      RECT 1.4520 0.6520 1.5020 0.8410 ;
      RECT 0.2050 0.5260 0.2550 0.8410 ;
      RECT 0.2790 0.8910 0.3290 1.2140 ;
      RECT 0.2050 0.4760 0.3290 0.5260 ;
      RECT 0.2790 0.3160 0.3290 0.4760 ;
      RECT 3.1670 0.8540 4.0690 0.9040 ;
      RECT 3.1670 0.6130 3.2170 0.8540 ;
      RECT 3.1670 0.9040 3.2170 1.0590 ;
      RECT 3.1670 0.5630 3.3690 0.6130 ;
      RECT 3.1670 1.0590 3.5370 1.1090 ;
      RECT 3.3190 0.4070 3.3690 0.5630 ;
      RECT 3.1670 0.4130 3.2170 0.5630 ;
      RECT 3.1670 1.1090 3.2170 1.3370 ;
      RECT 6.2830 0.6420 6.8050 0.6920 ;
      RECT 5.8180 0.4500 5.8680 0.7290 ;
      RECT 5.8180 0.7290 6.0050 0.7790 ;
      RECT 5.9550 0.7790 6.0050 1.1790 ;
      RECT 5.4480 1.1790 6.0050 1.2290 ;
      RECT 6.2830 0.4500 6.3330 0.6420 ;
      RECT 5.4470 0.4000 6.3330 0.4500 ;
      RECT 5.4470 0.4500 5.4970 0.5630 ;
      RECT 5.4470 0.2970 5.4970 0.4000 ;
      RECT 5.4480 1.2290 5.4980 1.3530 ;
      RECT 5.0310 0.5380 5.0810 1.0200 ;
      RECT 4.5190 0.5070 5.0810 0.5380 ;
      RECT 4.5350 1.0200 5.0810 1.0700 ;
      RECT 4.5190 0.4880 5.0800 0.5070 ;
      RECT 4.2710 0.7880 4.3210 1.1200 ;
      RECT 3.3740 0.7380 4.3230 0.7880 ;
      RECT 4.0790 0.5050 4.1290 0.7380 ;
      RECT 4.5350 1.0700 4.5850 1.1200 ;
      RECT 4.0580 1.1200 4.5850 1.1700 ;
      RECT 4.9950 0.1880 5.5890 0.2380 ;
      RECT 4.9950 0.2380 5.0450 0.2880 ;
      RECT 4.3540 0.2880 5.0450 0.3380 ;
      RECT 3.9470 0.4550 3.9970 0.6130 ;
      RECT 3.6830 0.6130 3.9970 0.6630 ;
      RECT 4.3540 0.3380 4.4040 0.4050 ;
      RECT 3.9470 0.4050 4.4040 0.4550 ;
      RECT 6.8700 0.6130 7.4130 0.6630 ;
      RECT 6.8700 0.6630 6.9200 0.7420 ;
      RECT 6.0550 0.7420 6.9200 0.7920 ;
      RECT 6.0550 0.7920 6.1050 1.3010 ;
      RECT 6.0550 0.6780 6.1050 0.7420 ;
      RECT 5.9630 0.6280 6.1050 0.6780 ;
      RECT 6.0550 0.5000 6.1050 0.6280 ;
      RECT 6.3590 0.7920 6.4090 1.3010 ;
      RECT 3.0150 0.8130 3.1050 0.8630 ;
      RECT 3.0550 0.4620 3.1050 0.8130 ;
      RECT 3.0150 0.8630 3.0650 1.0830 ;
      RECT 2.9990 0.4120 3.1050 0.4620 ;
      RECT 2.2550 1.0830 3.0650 1.1330 ;
      RECT 3.0150 1.1330 3.0650 1.3540 ;
      RECT 2.2550 0.7520 2.3050 1.0830 ;
      RECT 2.2550 0.7020 2.3450 0.7520 ;
      RECT 2.2950 0.5510 2.3450 0.7020 ;
      RECT 2.2550 0.5010 2.3450 0.5510 ;
      RECT 2.2550 0.4070 2.3050 0.5010 ;
      RECT 2.4070 0.6130 2.8530 0.6630 ;
      RECT 2.4070 0.6630 2.4570 1.0040 ;
      RECT 2.4070 0.4130 2.4570 0.6130 ;
      RECT 2.6180 0.0940 3.3150 0.1440 ;
      RECT 8.3190 0.8200 8.8670 0.8700 ;
      RECT 1.6500 0.7020 1.9410 0.7280 ;
      RECT 1.6870 0.6780 1.9410 0.7020 ;
      RECT 1.3430 0.4600 1.3930 0.5020 ;
      RECT 1.0230 0.4100 1.3930 0.4600 ;
      RECT 1.0230 1.0200 1.7000 1.0700 ;
      RECT 1.6500 0.7520 1.7000 1.0200 ;
      RECT 1.6500 0.7280 1.7370 0.7520 ;
      RECT 1.6870 0.5520 1.7370 0.6780 ;
      RECT 1.3430 0.5020 1.7370 0.5520 ;
      RECT 0.8870 0.3100 1.5450 0.3600 ;
      RECT 1.4950 0.3600 1.5450 0.3920 ;
      RECT 0.8870 0.3600 0.9370 0.3920 ;
      RECT 5.5070 0.8660 5.6560 0.9160 ;
      RECT 5.6060 0.9160 5.6560 0.9670 ;
      RECT 5.6060 0.9670 5.7410 1.0170 ;
      RECT 1.9910 0.6280 2.2450 0.6520 ;
      RECT 1.9520 0.6020 2.2450 0.6280 ;
      RECT 1.9910 0.6520 2.0410 0.7780 ;
      RECT 1.9520 0.5780 2.0410 0.6020 ;
      RECT 1.9520 0.7780 2.0410 0.8280 ;
      RECT 1.9520 0.3190 2.0020 0.5780 ;
      RECT 1.9520 0.8280 2.0020 1.0760 ;
      RECT 8.6230 0.7090 9.1610 0.7590 ;
      RECT 7.8790 1.0920 8.3280 1.1420 ;
      RECT 7.8790 0.6770 7.9290 1.0920 ;
      RECT 7.8390 0.6270 7.9290 0.6770 ;
      RECT 7.8390 0.4770 7.8890 0.6270 ;
      RECT 7.8390 0.4270 7.9290 0.4770 ;
      RECT 7.8790 0.1260 7.9290 0.4270 ;
      RECT 8.8510 1.0950 9.3890 1.1450 ;
      RECT 8.3190 0.2480 9.1610 0.2980 ;
      RECT 5.0490 1.5200 8.3250 1.5700 ;
      RECT 9.2470 0.6770 9.2970 0.7680 ;
      RECT 9.2070 0.4270 9.2970 0.4620 ;
      RECT 9.2470 0.1260 9.2970 0.4270 ;
      RECT 9.2070 0.6270 9.2970 0.6770 ;
      RECT 9.2070 0.5120 9.2570 0.6270 ;
      RECT 9.0030 0.4770 9.2570 0.5120 ;
      RECT 9.0030 0.4620 9.2970 0.4770 ;
      RECT 4.2910 1.5200 4.9810 1.5700 ;
      RECT 4.7460 0.6130 4.9810 0.6630 ;
      RECT 5.2950 0.8670 5.4370 0.9170 ;
      RECT 5.2950 0.6630 5.3450 0.8670 ;
      RECT 5.2950 0.6130 5.7410 0.6630 ;
      RECT 4.3830 0.9200 4.8130 0.9700 ;
      RECT 4.7630 0.8310 4.8130 0.9200 ;
      RECT 4.3830 0.9700 4.4330 1.0340 ;
      RECT 4.3830 0.5050 4.4330 0.9200 ;
      RECT 4.1390 1.4200 5.4450 1.4700 ;
      RECT 3.3030 1.1900 3.6890 1.2400 ;
      RECT 3.2270 1.3890 3.7650 1.4390 ;
      RECT 7.3310 1.2340 8.6290 1.2840 ;
      RECT 7.9390 0.5270 8.5370 0.5770 ;
      RECT 8.4870 0.5770 8.5370 0.7700 ;
      RECT 8.4870 0.3480 8.5370 0.5270 ;
      RECT 8.1830 0.5770 8.2330 0.8870 ;
      RECT 8.1830 0.1260 8.2330 0.5270 ;
      RECT 8.6230 0.1320 8.8570 0.1820 ;
      RECT 2.9230 1.5240 3.9170 1.5740 ;
      RECT 5.8110 0.0940 6.0450 0.1440 ;
      RECT 0.7190 0.5100 1.2570 0.5600 ;
      RECT 1.1750 1.1330 1.5610 1.1830 ;
      RECT 0.7190 0.9410 0.9530 0.9910 ;
      RECT 2.8630 0.7130 2.9890 0.7630 ;
      RECT 2.8630 0.7630 2.9130 1.0330 ;
      RECT 2.9390 0.5630 2.9890 0.7130 ;
      RECT 2.8470 0.5130 2.9890 0.5630 ;
      RECT 4.6710 0.3880 5.3450 0.4380 ;
      RECT 5.2950 0.4380 5.3450 0.5630 ;
      RECT 5.2950 0.2970 5.3450 0.3880 ;
      RECT 5.1430 0.3840 5.1930 0.3880 ;
      RECT 5.1430 0.4380 5.1930 0.9670 ;
      RECT 5.1430 0.9670 5.3610 1.0170 ;
    LAYER PO ;
      RECT 7.3570 0.0670 7.3870 1.6050 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 4.9250 0.8390 4.9550 1.6060 ;
      RECT 9.4850 0.0660 9.5150 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 5.6850 0.0660 5.7150 0.6910 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 3.1010 0.8400 3.1310 1.6060 ;
      RECT 5.6850 0.9390 5.7150 1.6060 ;
      RECT 5.3810 0.0660 5.4110 0.6370 ;
      RECT 3.1010 0.0660 3.1310 0.6370 ;
      RECT 3.7090 0.0660 3.7390 0.6910 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 9.3330 0.0660 9.3630 1.6060 ;
      RECT 4.9250 0.0660 4.9550 0.6910 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 9.6370 0.0660 9.6670 1.6060 ;
      RECT 4.6210 0.8920 4.6510 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 5.3810 0.8390 5.4110 1.6060 ;
      RECT 9.7890 0.0660 9.8190 1.6060 ;
      RECT 10.2450 0.0660 10.2750 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 9.9410 0.0660 9.9710 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 10.0930 0.0660 10.1230 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 4.6210 0.0660 4.6510 0.6910 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 3.7090 0.9390 3.7390 1.6060 ;
    LAYER NWELL ;
      RECT 7.7120 0.4910 9.7230 1.0830 ;
      RECT -0.1150 1.5430 10.4580 1.7730 ;
      RECT -0.1150 0.6790 7.2500 1.5430 ;
      RECT 10.1830 0.6790 10.4580 1.5430 ;
  END
END RSDFFSRARX2_LVT

MACRO RDFFSRSSRX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.12 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 9.1200 1.7020 ;
        RECT 1.1910 1.1310 1.2410 1.6420 ;
        RECT 0.2790 1.3460 0.3290 1.6420 ;
        RECT 1.7990 1.3880 1.8490 1.6420 ;
        RECT 3.0550 1.2700 3.1050 1.6420 ;
        RECT 7.1590 1.4540 7.2090 1.6420 ;
        RECT 0.2790 1.2960 0.6330 1.3460 ;
        RECT 1.6270 1.3380 1.8490 1.3880 ;
        RECT 2.8460 1.2200 3.9930 1.2700 ;
        RECT 4.6870 1.4040 7.2090 1.4540 ;
        RECT 0.2790 0.9300 0.3290 1.2960 ;
        RECT 0.5830 0.9800 0.6330 1.2960 ;
        RECT 4.6870 1.2790 4.7370 1.4040 ;
        RECT 5.7510 0.9590 5.8010 1.4040 ;
        RECT 5.2950 0.9530 5.3450 1.4040 ;
    END
  END VDD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.5990 0.4010 6.2990 0.4510 ;
        RECT 5.5990 0.1570 5.6490 0.4010 ;
        RECT 6.1770 0.4510 6.2990 0.5380 ;
        RECT 6.2490 0.5380 6.2990 0.8590 ;
        RECT 5.5990 0.8590 6.2990 0.9090 ;
        RECT 5.5990 0.9090 5.6490 1.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.9030 0.9690 6.4370 1.0190 ;
        RECT 6.3870 0.3510 6.4370 0.9690 ;
        RECT 5.9030 1.0190 6.1350 1.1290 ;
        RECT 5.8870 0.3010 6.4370 0.3510 ;
        RECT 5.9030 1.1290 5.9530 1.3270 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.5550 1.4650 1.7270 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 9.1200 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.3550 ;
        RECT 1.5710 0.0300 1.6210 0.2740 ;
        RECT 8.1830 0.0300 8.2330 0.4260 ;
        RECT 5.7510 0.0300 5.8010 0.2410 ;
        RECT 6.8150 0.0300 6.8650 0.4260 ;
        RECT 1.1910 0.0300 1.2410 0.4050 ;
        RECT 7.7270 0.0300 7.7770 0.1980 ;
        RECT 5.4710 0.0300 5.5210 0.3000 ;
        RECT 0.2790 0.3550 0.6330 0.4050 ;
        RECT 1.5710 0.2740 3.0650 0.3240 ;
        RECT 4.6710 0.3000 5.5210 0.3500 ;
        RECT 0.5830 0.4050 0.6330 0.5290 ;
        RECT 0.2790 0.4050 0.3290 0.5130 ;
        RECT 3.0150 0.3240 3.0650 0.3470 ;
        RECT 2.8630 0.3240 2.9130 0.5570 ;
        RECT 1.6470 0.3240 1.6970 0.5570 ;
        RECT 1.7990 0.3240 1.8490 0.5570 ;
        RECT 3.0150 0.2470 3.0650 0.2740 ;
        RECT 3.0150 0.1970 3.9930 0.2470 ;
        RECT 3.3190 0.2470 3.3690 0.3490 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9470 0.8570 1.1190 0.9770 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7010 0.4210 0.7510 ;
        RECT 0.2490 0.7510 0.3590 0.8250 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SETB

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.3050 0.2490 8.4170 0.3590 ;
        RECT 8.3160 0.3590 8.3660 0.5080 ;
        RECT 8.0910 0.5080 8.3660 0.5580 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.5930 0.7050 3.7490 0.7310 ;
        RECT 3.5930 0.7310 4.0530 0.7810 ;
        RECT 3.6990 0.5970 3.7490 0.7050 ;
        RECT 3.5930 0.7810 3.7490 0.8150 ;
        RECT 4.0030 0.7810 4.0530 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 0.0970 0.5110 0.1910 ;
        RECT 0.4010 0.1910 0.7250 0.2410 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END RSTB

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 6.7990 0.9420 8.4170 1.0020 ;
        RECT 8.3070 0.6900 8.4170 0.9420 ;
        RECT 8.1830 0.6270 8.2330 0.9420 ;
    END
  END VDDG
  OBS
    LAYER M1 ;
      RECT 4.9060 0.7290 5.0930 0.7790 ;
      RECT 5.0430 0.7790 5.0930 1.1790 ;
      RECT 4.5360 1.1790 5.0930 1.2290 ;
      RECT 5.3710 0.4500 5.4210 0.6580 ;
      RECT 4.5350 0.4000 5.4210 0.4500 ;
      RECT 4.5350 0.4500 4.5850 0.5630 ;
      RECT 4.5350 0.2970 4.5850 0.4000 ;
      RECT 4.5360 1.2290 4.5860 1.3530 ;
      RECT 4.5950 0.8660 4.7440 0.9160 ;
      RECT 4.6940 0.9160 4.7440 0.9670 ;
      RECT 4.6940 0.9670 4.8290 1.0170 ;
      RECT 5.2190 0.0920 5.2690 0.2000 ;
      RECT 4.7270 0.2000 5.2690 0.2500 ;
      RECT 4.7270 0.1470 4.7770 0.2000 ;
      RECT 2.6190 0.0970 4.7770 0.1470 ;
      RECT 5.7750 0.6130 6.1970 0.6630 ;
      RECT 5.1430 0.8090 5.1930 1.3010 ;
      RECT 5.1430 0.6780 5.1930 0.7590 ;
      RECT 5.0510 0.6280 5.1930 0.6780 ;
      RECT 5.1430 0.5000 5.1930 0.6280 ;
      RECT 5.4470 0.8090 5.4970 1.3010 ;
      RECT 5.7750 0.6630 5.8250 0.7590 ;
      RECT 5.1430 0.7590 5.8250 0.8090 ;
      RECT 2.1030 0.8130 2.1930 0.8630 ;
      RECT 2.1430 0.4620 2.1930 0.8130 ;
      RECT 2.1030 0.8630 2.1530 1.2020 ;
      RECT 2.0870 0.4120 2.1930 0.4620 ;
      RECT 1.3430 1.2020 2.1530 1.2520 ;
      RECT 2.1030 1.2520 2.1530 1.3540 ;
      RECT 1.3430 0.8690 1.3930 1.2020 ;
      RECT 1.3430 0.8190 1.4330 0.8690 ;
      RECT 1.3830 0.4750 1.4330 0.8190 ;
      RECT 1.3430 0.4250 1.4330 0.4750 ;
      RECT 1.3430 0.3620 1.3930 0.4250 ;
      RECT 7.4070 0.7090 7.9450 0.7590 ;
      RECT 0.7350 1.3160 1.1060 1.3660 ;
      RECT 0.7350 0.9800 0.7850 1.3160 ;
      RECT 1.4950 0.6130 1.9410 0.6630 ;
      RECT 1.4950 0.6630 1.5450 1.0040 ;
      RECT 1.4950 0.4130 1.5450 0.6130 ;
      RECT 4.1190 0.5470 4.1690 1.0200 ;
      RECT 3.6230 1.0200 4.1690 1.0700 ;
      RECT 3.6070 0.4970 4.1680 0.5070 ;
      RECT 3.6070 0.5070 4.1690 0.5470 ;
      RECT 3.3590 0.7880 3.4090 1.1200 ;
      RECT 2.4620 0.7380 3.4110 0.7880 ;
      RECT 3.1670 0.5050 3.2170 0.7380 ;
      RECT 3.6230 1.0700 3.6730 1.1200 ;
      RECT 3.1460 1.1200 3.6730 1.1700 ;
      RECT 7.9910 0.6270 8.0810 0.6770 ;
      RECT 8.0310 0.6770 8.0810 0.7680 ;
      RECT 7.9910 0.3980 8.0810 0.4480 ;
      RECT 8.0310 0.1260 8.0810 0.3980 ;
      RECT 7.9910 0.5120 8.0410 0.6270 ;
      RECT 7.7870 0.4620 8.0410 0.5120 ;
      RECT 7.9910 0.4480 8.0410 0.4620 ;
      RECT 3.3790 1.5200 4.0690 1.5700 ;
      RECT 3.8340 0.6310 4.0690 0.6810 ;
      RECT 4.3830 0.8670 4.5250 0.9170 ;
      RECT 4.3830 0.7220 4.4330 0.8670 ;
      RECT 4.3830 0.6720 4.8290 0.7220 ;
      RECT 3.4710 0.9200 3.9010 0.9700 ;
      RECT 3.8510 0.8310 3.9010 0.9200 ;
      RECT 3.4710 0.9700 3.5210 1.0340 ;
      RECT 3.4710 0.5050 3.5210 0.9200 ;
      RECT 3.2270 1.4200 4.5330 1.4700 ;
      RECT 2.3910 1.1900 2.7770 1.2400 ;
      RECT 2.3150 1.3890 2.8530 1.4390 ;
      RECT 4.0830 0.1970 4.6770 0.2470 ;
      RECT 4.0830 0.2470 4.1330 0.2970 ;
      RECT 3.4420 0.2970 4.1330 0.3470 ;
      RECT 3.0350 0.4550 3.0850 0.6130 ;
      RECT 2.7710 0.6130 3.0850 0.6630 ;
      RECT 3.4420 0.3470 3.4920 0.4050 ;
      RECT 3.0350 0.4050 3.4920 0.4550 ;
      RECT 0.9560 0.6240 1.3330 0.6740 ;
      RECT 0.9560 0.4930 1.0060 0.6240 ;
      RECT 0.9560 0.6740 1.0060 0.7520 ;
      RECT 0.8710 0.4430 1.0060 0.4930 ;
      RECT 0.8470 0.7520 1.0060 0.8020 ;
      RECT 0.8470 1.0470 0.9370 1.0970 ;
      RECT 0.8870 1.0970 0.9370 1.2460 ;
      RECT 0.8470 0.8020 0.8970 1.0470 ;
      RECT 6.1150 1.1990 7.4130 1.2490 ;
      RECT 1.7060 0.0940 2.4030 0.1440 ;
      RECT 7.1030 0.8200 7.6510 0.8700 ;
      RECT 0.7000 0.5730 0.8770 0.6230 ;
      RECT 0.7000 0.6230 0.7500 0.8440 ;
      RECT 0.4310 0.8440 0.7500 0.8940 ;
      RECT 0.4310 0.8940 0.4810 1.2460 ;
      RECT 0.4310 0.4550 0.4810 0.6010 ;
      RECT 0.4710 0.6510 0.5210 0.8440 ;
      RECT 0.4310 0.6010 0.5210 0.6510 ;
      RECT 7.4070 0.1320 7.6410 0.1820 ;
      RECT 6.6630 1.0740 7.1120 1.1240 ;
      RECT 6.6630 0.6770 6.7130 1.0740 ;
      RECT 6.6230 0.6270 6.7130 0.6770 ;
      RECT 6.6230 0.4770 6.6730 0.6270 ;
      RECT 6.6230 0.4270 6.7130 0.4770 ;
      RECT 6.6630 0.1260 6.7130 0.4270 ;
      RECT 0.7190 0.3010 1.1050 0.3510 ;
      RECT 2.0110 1.5240 3.0050 1.5740 ;
      RECT 6.7230 0.5270 7.3210 0.5770 ;
      RECT 6.9670 0.5770 7.0170 0.8690 ;
      RECT 6.9670 0.1260 7.0170 0.5270 ;
      RECT 7.2710 0.5770 7.3210 0.7700 ;
      RECT 7.2710 0.3480 7.3210 0.5270 ;
      RECT 0.4910 1.4490 0.8770 1.4990 ;
      RECT 4.8990 0.0940 5.1330 0.1440 ;
      RECT 7.6350 1.0770 8.1730 1.1270 ;
      RECT 7.1030 0.2480 7.9450 0.2980 ;
      RECT 4.1370 1.5200 7.1090 1.5700 ;
      RECT 1.9510 0.7130 2.0770 0.7630 ;
      RECT 1.9510 0.7630 2.0010 1.0330 ;
      RECT 2.0270 0.5630 2.0770 0.7130 ;
      RECT 1.9350 0.5130 2.0770 0.5630 ;
      RECT 3.7590 0.3970 4.4330 0.4470 ;
      RECT 4.3830 0.4470 4.4330 0.5630 ;
      RECT 4.3830 0.2970 4.4330 0.3970 ;
      RECT 4.2310 0.4470 4.2810 0.9670 ;
      RECT 4.2310 0.9670 4.4490 1.0170 ;
      RECT 4.2310 1.0170 4.2810 1.1200 ;
      RECT 4.2310 1.1700 4.2810 1.2700 ;
      RECT 3.7590 1.1200 4.2810 1.1700 ;
      RECT 3.2090 0.8580 3.3090 0.9080 ;
      RECT 3.2090 0.9080 3.2590 0.9680 ;
      RECT 2.7710 0.9680 3.2590 1.0180 ;
      RECT 2.2550 0.8540 3.1570 0.9040 ;
      RECT 2.2550 0.9040 2.3050 1.0590 ;
      RECT 2.2550 0.6130 2.3050 0.8540 ;
      RECT 2.2550 1.0590 2.6250 1.1090 ;
      RECT 2.2550 0.5630 2.4570 0.6130 ;
      RECT 2.2550 1.1090 2.3050 1.3370 ;
      RECT 2.4070 0.4070 2.4570 0.5630 ;
      RECT 2.2550 0.4130 2.3050 0.5630 ;
      RECT 5.3710 0.6580 5.7250 0.7080 ;
      RECT 5.6750 0.6230 5.7250 0.6580 ;
      RECT 4.9060 0.4500 4.9560 0.7290 ;
    LAYER PO ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 2.1890 0.8400 2.2190 1.6060 ;
      RECT 4.7730 0.9390 4.8030 1.6060 ;
      RECT 4.4690 0.0660 4.4990 0.6550 ;
      RECT 2.1890 0.0660 2.2190 0.6370 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 2.7970 0.0660 2.8270 0.6910 ;
      RECT 4.0130 0.0660 4.0430 0.6910 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 0.6690 0.0760 0.6990 0.5970 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 3.7090 0.8920 3.7390 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 4.4690 0.8390 4.4990 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 0.8210 0.8700 0.8510 1.6060 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 0.5170 0.0760 0.5470 1.6060 ;
      RECT 0.8210 0.0760 0.8510 0.6510 ;
      RECT 0.6690 0.8160 0.6990 1.6060 ;
      RECT 0.3650 0.0760 0.3950 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 3.7090 0.0660 3.7390 0.6910 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 2.7970 0.9390 2.8270 1.6060 ;
      RECT 6.1410 0.0670 6.1710 1.6050 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 4.0130 0.8390 4.0430 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 4.7730 0.0660 4.8030 0.7540 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
    LAYER NWELL ;
      RECT 6.4960 0.4910 8.5070 1.0830 ;
      RECT -0.1150 1.5430 9.2410 1.7730 ;
      RECT -0.1150 0.6790 6.0340 1.5430 ;
      RECT 8.9670 0.6790 9.2410 1.5430 ;
  END
END RDFFSRSSRX1_LVT

MACRO RDFFSRSSRX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.424 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.6330 0.3210 6.7530 0.3600 ;
        RECT 6.0550 0.2710 6.7530 0.3210 ;
        RECT 6.7030 0.3600 6.7530 0.9330 ;
        RECT 6.6330 0.2500 6.7530 0.2710 ;
        RECT 6.0550 0.1490 6.1050 0.2710 ;
        RECT 6.0550 0.9330 6.7530 0.9830 ;
        RECT 6.6330 0.2490 6.7450 0.2500 ;
        RECT 6.0550 0.9830 6.1050 1.3270 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 9.4240 1.7020 ;
        RECT 1.1910 1.1310 1.2410 1.6420 ;
        RECT 7.4630 1.4540 7.5130 1.6420 ;
        RECT 0.2790 1.3460 0.3290 1.6420 ;
        RECT 1.7990 1.3880 1.8490 1.6420 ;
        RECT 3.0550 1.2700 3.1050 1.6420 ;
        RECT 4.6870 1.4040 7.5130 1.4540 ;
        RECT 0.2790 1.2960 0.6330 1.3460 ;
        RECT 1.6270 1.3380 1.8490 1.3880 ;
        RECT 2.8460 1.2200 3.9930 1.2700 ;
        RECT 4.6870 1.2790 4.7370 1.4040 ;
        RECT 5.9030 0.9610 5.9530 1.4040 ;
        RECT 5.5990 0.9130 5.6490 1.4040 ;
        RECT 5.2950 0.9530 5.3450 1.4040 ;
        RECT 6.2070 1.0530 6.2570 1.4040 ;
        RECT 0.2790 0.9300 0.3290 1.2960 ;
        RECT 0.5830 0.9800 0.6330 1.2960 ;
    END
  END VDD

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.5550 1.4650 1.7270 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 9.4240 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.3550 ;
        RECT 1.5710 0.0300 1.6210 0.2740 ;
        RECT 8.4870 0.0300 8.5370 0.4260 ;
        RECT 5.5990 0.0300 5.6490 0.4090 ;
        RECT 6.2070 0.0300 6.2570 0.2210 ;
        RECT 5.9030 0.0300 5.9530 0.3200 ;
        RECT 7.1190 0.0300 7.1690 0.4260 ;
        RECT 1.1910 0.0300 1.2410 0.4050 ;
        RECT 8.0310 0.0300 8.0810 0.1980 ;
        RECT 5.4710 0.0300 5.5210 0.3000 ;
        RECT 0.2790 0.3550 0.6330 0.4050 ;
        RECT 1.5710 0.2740 3.0650 0.3240 ;
        RECT 4.6710 0.3000 5.5210 0.3500 ;
        RECT 0.5830 0.4050 0.6330 0.5290 ;
        RECT 0.2790 0.4050 0.3290 0.5130 ;
        RECT 3.0150 0.3240 3.0650 0.3470 ;
        RECT 2.8630 0.3240 2.9130 0.5570 ;
        RECT 1.6470 0.3240 1.6970 0.5570 ;
        RECT 1.7990 0.3240 1.8490 0.5570 ;
        RECT 3.0150 0.2380 3.0650 0.2740 ;
        RECT 3.0150 0.1880 3.9930 0.2380 ;
        RECT 3.3190 0.2380 3.3690 0.3490 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9470 0.8570 1.1190 0.9770 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7010 0.4210 0.7510 ;
        RECT 0.2490 0.7510 0.3590 0.8250 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SETB

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.6090 0.2490 8.7210 0.3590 ;
        RECT 8.6200 0.3590 8.6700 0.5270 ;
        RECT 8.3950 0.5270 8.6700 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.5930 0.7050 3.7490 0.7310 ;
        RECT 3.5930 0.7310 4.0530 0.7810 ;
        RECT 3.6990 0.5970 3.7490 0.7050 ;
        RECT 3.5930 0.7810 3.7490 0.8150 ;
        RECT 4.0030 0.7810 4.0530 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 0.0970 0.5110 0.1910 ;
        RECT 0.4010 0.1910 0.7250 0.2410 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END RSTB

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.4810 0.4010 6.5930 0.4020 ;
        RECT 5.7510 0.4020 6.6030 0.4520 ;
        RECT 5.7510 0.1490 5.8010 0.4020 ;
        RECT 6.4810 0.4520 6.6030 0.5120 ;
        RECT 6.5530 0.5120 6.6030 0.8330 ;
        RECT 5.7510 0.8330 6.6030 0.8830 ;
        RECT 5.7510 0.8830 5.8010 1.3190 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 7.1030 0.9420 8.7210 1.0020 ;
        RECT 8.6110 0.6900 8.7210 0.9420 ;
        RECT 8.4870 0.6270 8.5370 0.9420 ;
    END
  END VDDG
  OBS
    LAYER M1 ;
      RECT 4.9060 0.4500 4.9560 0.7290 ;
      RECT 4.9060 0.7290 5.0930 0.7790 ;
      RECT 5.0430 0.7790 5.0930 1.1790 ;
      RECT 4.5360 1.1790 5.0930 1.2290 ;
      RECT 5.3710 0.4500 5.4210 0.6320 ;
      RECT 4.5350 0.4000 5.4210 0.4500 ;
      RECT 0.9560 0.6240 1.3330 0.6740 ;
      RECT 0.9560 0.4930 1.0060 0.6240 ;
      RECT 0.9560 0.6740 1.0060 0.7520 ;
      RECT 0.8710 0.4430 1.0060 0.4930 ;
      RECT 0.8470 0.7520 1.0060 0.8020 ;
      RECT 0.8470 1.0470 0.9370 1.0970 ;
      RECT 0.8870 1.0970 0.9370 1.2460 ;
      RECT 0.8470 0.8020 0.8970 1.0470 ;
      RECT 0.7000 0.5730 0.8770 0.6230 ;
      RECT 0.7000 0.6230 0.7500 0.8440 ;
      RECT 0.4310 0.8440 0.7500 0.8940 ;
      RECT 0.4310 0.8940 0.4810 1.2460 ;
      RECT 0.4310 0.4550 0.4810 0.6010 ;
      RECT 0.4710 0.6510 0.5210 0.8440 ;
      RECT 0.4310 0.6010 0.5210 0.6510 ;
      RECT 4.5950 0.8660 4.7440 0.9160 ;
      RECT 4.6940 0.9160 4.7440 0.9670 ;
      RECT 4.6940 0.9670 4.8290 1.0170 ;
      RECT 4.7270 0.2000 5.2690 0.2500 ;
      RECT 5.2190 0.0880 5.2690 0.2000 ;
      RECT 4.7270 0.1380 4.7770 0.2000 ;
      RECT 2.6190 0.0880 4.7770 0.1380 ;
      RECT 5.9430 0.6130 6.5010 0.6630 ;
      RECT 5.1430 0.7820 5.1930 1.3010 ;
      RECT 5.1430 0.6780 5.1930 0.7320 ;
      RECT 5.0510 0.6280 5.1930 0.6780 ;
      RECT 5.1430 0.5000 5.1930 0.6280 ;
      RECT 5.4470 0.7820 5.4970 1.3010 ;
      RECT 5.9430 0.6630 5.9930 0.7320 ;
      RECT 5.1430 0.7320 5.9930 0.7820 ;
      RECT 2.1030 0.8130 2.1930 0.8630 ;
      RECT 2.1430 0.4620 2.1930 0.8130 ;
      RECT 2.1030 0.8630 2.1530 1.2020 ;
      RECT 2.0870 0.4120 2.1930 0.4620 ;
      RECT 1.3430 1.2020 2.1530 1.2520 ;
      RECT 2.1030 1.2520 2.1530 1.3540 ;
      RECT 1.3430 0.8690 1.3930 1.2020 ;
      RECT 1.3430 0.8190 1.4330 0.8690 ;
      RECT 1.3830 0.4750 1.4330 0.8190 ;
      RECT 1.3430 0.4250 1.4330 0.4750 ;
      RECT 1.3430 0.3620 1.3930 0.4250 ;
      RECT 7.7110 0.7090 8.2490 0.7590 ;
      RECT 0.7350 1.3160 1.1060 1.3660 ;
      RECT 0.7350 0.9800 0.7850 1.3160 ;
      RECT 3.6070 0.4880 4.1680 0.5110 ;
      RECT 3.6070 0.5110 4.1690 0.5380 ;
      RECT 4.1190 0.5380 4.1690 1.0200 ;
      RECT 3.6230 1.0200 4.1690 1.0700 ;
      RECT 3.3590 0.7880 3.4090 1.1200 ;
      RECT 2.4620 0.7380 3.4110 0.7880 ;
      RECT 3.1670 0.5050 3.2170 0.7380 ;
      RECT 3.6230 1.0700 3.6730 1.1200 ;
      RECT 3.1460 1.1200 3.6730 1.1700 ;
      RECT 4.1370 1.5200 7.4130 1.5700 ;
      RECT 1.4950 0.6130 1.9410 0.6630 ;
      RECT 1.4950 0.6630 1.5450 1.0040 ;
      RECT 1.4950 0.4130 1.5450 0.6130 ;
      RECT 8.3350 0.6770 8.3850 0.7680 ;
      RECT 8.2950 0.4270 8.3850 0.4620 ;
      RECT 8.3350 0.1260 8.3850 0.4270 ;
      RECT 8.2950 0.6270 8.3850 0.6770 ;
      RECT 8.2950 0.5120 8.3450 0.6270 ;
      RECT 8.0910 0.4770 8.3450 0.5120 ;
      RECT 8.0910 0.4620 8.3850 0.4770 ;
      RECT 3.3790 1.5200 4.0690 1.5700 ;
      RECT 3.8340 0.6130 4.0690 0.6630 ;
      RECT 4.3830 0.8670 4.5250 0.9170 ;
      RECT 4.3830 0.6630 4.4330 0.8670 ;
      RECT 4.3830 0.6130 4.8290 0.6630 ;
      RECT 3.4710 0.9200 3.9010 0.9700 ;
      RECT 3.8510 0.8310 3.9010 0.9200 ;
      RECT 3.4710 0.9700 3.5210 1.0340 ;
      RECT 3.4710 0.5050 3.5210 0.9200 ;
      RECT 3.2270 1.4200 4.5330 1.4700 ;
      RECT 2.3910 1.1900 2.7770 1.2400 ;
      RECT 2.3150 1.3890 2.8530 1.4390 ;
      RECT 4.0830 0.1880 4.6770 0.2380 ;
      RECT 4.0830 0.2380 4.1330 0.2880 ;
      RECT 3.4420 0.2880 4.1330 0.3380 ;
      RECT 3.0350 0.4550 3.0850 0.6130 ;
      RECT 2.7710 0.6130 3.0850 0.6630 ;
      RECT 3.4420 0.3380 3.4920 0.4050 ;
      RECT 3.0350 0.4050 3.4920 0.4550 ;
      RECT 6.4190 1.1990 7.7170 1.2490 ;
      RECT 1.7060 0.0940 2.4030 0.1440 ;
      RECT 7.4070 0.8200 7.9550 0.8700 ;
      RECT 7.7110 0.1320 7.9450 0.1820 ;
      RECT 6.9670 1.0620 7.4160 1.1120 ;
      RECT 6.9670 0.6770 7.0170 1.0620 ;
      RECT 6.9270 0.6270 7.0170 0.6770 ;
      RECT 6.9270 0.4770 6.9770 0.6270 ;
      RECT 6.9270 0.4270 7.0170 0.4770 ;
      RECT 6.9670 0.1260 7.0170 0.4270 ;
      RECT 0.7190 0.3010 1.1050 0.3510 ;
      RECT 2.0110 1.5240 3.0050 1.5740 ;
      RECT 7.0270 0.5270 7.6250 0.5770 ;
      RECT 7.2710 0.5770 7.3210 0.8840 ;
      RECT 7.2710 0.1260 7.3210 0.5270 ;
      RECT 7.5750 0.5770 7.6250 0.7700 ;
      RECT 7.5750 0.3480 7.6250 0.5270 ;
      RECT 0.4910 1.4490 0.8770 1.4990 ;
      RECT 4.8990 0.0940 5.1330 0.1440 ;
      RECT 7.9390 1.0620 8.4770 1.1120 ;
      RECT 7.4070 0.2480 8.2490 0.2980 ;
      RECT 1.9510 0.7130 2.0770 0.7630 ;
      RECT 1.9510 0.7630 2.0010 1.0330 ;
      RECT 2.0270 0.5630 2.0770 0.7130 ;
      RECT 1.9350 0.5130 2.0770 0.5630 ;
      RECT 3.7590 0.3880 4.4330 0.4380 ;
      RECT 4.3830 0.4380 4.4330 0.5630 ;
      RECT 4.3830 0.2970 4.4330 0.3880 ;
      RECT 4.2310 0.4380 4.2810 0.9670 ;
      RECT 4.2310 0.9670 4.4490 1.0170 ;
      RECT 4.2310 1.0170 4.2810 1.1200 ;
      RECT 4.2310 1.1700 4.2810 1.2700 ;
      RECT 3.7590 1.1200 4.2810 1.1700 ;
      RECT 3.2090 0.8580 3.3090 0.9080 ;
      RECT 3.2090 0.9080 3.2590 0.9680 ;
      RECT 2.7710 0.9680 3.2590 1.0180 ;
      RECT 2.2550 0.8540 3.1570 0.9040 ;
      RECT 2.2550 0.6130 2.3050 0.8540 ;
      RECT 2.2550 0.9040 2.3050 1.0590 ;
      RECT 2.2550 0.5630 2.4570 0.6130 ;
      RECT 2.2550 1.0590 2.6250 1.1090 ;
      RECT 2.4070 0.4070 2.4570 0.5630 ;
      RECT 2.2550 0.4130 2.3050 0.5630 ;
      RECT 2.2550 1.1090 2.3050 1.3370 ;
      RECT 5.3330 0.6320 5.8930 0.6820 ;
      RECT 4.5350 0.4500 4.5850 0.5630 ;
      RECT 4.5350 0.2970 4.5850 0.4000 ;
      RECT 4.5360 1.2290 4.5860 1.3530 ;
    LAYER PO ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 2.1890 0.8400 2.2190 1.6060 ;
      RECT 4.7730 0.9390 4.8030 1.6060 ;
      RECT 4.4690 0.0660 4.4990 0.6370 ;
      RECT 2.1890 0.0660 2.2190 0.6370 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 2.7970 0.0660 2.8270 0.6910 ;
      RECT 4.0130 0.0660 4.0430 0.6910 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 0.6690 0.0760 0.6990 0.5970 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 3.7090 0.8920 3.7390 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 4.4690 0.8390 4.4990 1.6060 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 9.3330 0.0660 9.3630 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 0.8210 0.8700 0.8510 1.6060 ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 0.5170 0.0760 0.5470 1.6060 ;
      RECT 0.8210 0.0760 0.8510 0.6510 ;
      RECT 0.6690 0.8160 0.6990 1.6060 ;
      RECT 0.3650 0.0760 0.3950 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 3.7090 0.0660 3.7390 0.6910 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 2.7970 0.9390 2.8270 1.6060 ;
      RECT 6.4450 0.0670 6.4750 1.6050 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 4.0130 0.8390 4.0430 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 4.7730 0.0660 4.8030 0.6910 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
    LAYER NWELL ;
      RECT 6.8000 0.4910 8.8110 1.0830 ;
      RECT -0.1150 1.5430 9.5460 1.7730 ;
      RECT -0.1150 0.6790 6.3380 1.5430 ;
      RECT 9.2710 0.6790 9.5460 1.5430 ;
  END
END RDFFSRSSRX2_LVT

MACRO RDFFSRX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.904 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 7.9040 1.7020 ;
        RECT 0.2790 1.1310 0.3290 1.6420 ;
        RECT 1.9910 1.2700 2.0410 1.6420 ;
        RECT 5.9430 1.4540 5.9930 1.6420 ;
        RECT 0.8870 1.2940 0.9370 1.6420 ;
        RECT 1.7830 1.2200 2.9290 1.2700 ;
        RECT 3.6230 1.4040 5.9930 1.4540 ;
        RECT 0.7150 1.2440 0.9370 1.2940 ;
        RECT 3.6230 1.2790 3.6730 1.4040 ;
        RECT 4.5350 0.9590 4.5850 1.4040 ;
        RECT 4.0790 0.9530 4.1290 1.4040 ;
    END
  END VDD

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.3830 0.4010 5.0830 0.4510 ;
        RECT 4.3830 0.1570 4.4330 0.4010 ;
        RECT 4.9610 0.4510 5.0830 0.5380 ;
        RECT 5.0330 0.5380 5.0830 0.8590 ;
        RECT 4.3830 0.8590 5.0830 0.9090 ;
        RECT 4.3830 0.9090 4.4330 1.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6870 0.9690 5.2210 1.0190 ;
        RECT 5.1710 0.3510 5.2210 0.9690 ;
        RECT 4.6870 1.0190 4.9190 1.1290 ;
        RECT 4.6710 0.3010 5.2210 0.3510 ;
        RECT 4.6870 1.1290 4.7370 1.3270 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6430 1.4650 0.8150 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 7.9040 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.2570 ;
        RECT 6.5110 0.0300 6.5610 0.1980 ;
        RECT 6.9670 0.0300 7.0170 0.4260 ;
        RECT 4.5350 0.0300 4.5850 0.2410 ;
        RECT 5.5990 0.0300 5.6490 0.4260 ;
        RECT 4.2550 0.0300 4.3050 0.2830 ;
        RECT 0.2790 0.2570 2.0010 0.3070 ;
        RECT 3.6070 0.2830 4.3050 0.3330 ;
        RECT 0.7350 0.3070 0.7850 0.5570 ;
        RECT 0.8870 0.3070 0.9370 0.5570 ;
        RECT 0.2790 0.3070 0.3290 0.4050 ;
        RECT 1.9510 0.2340 2.0010 0.2570 ;
        RECT 1.9510 0.1840 2.9290 0.2340 ;
        RECT 2.2550 0.2340 2.3050 0.3490 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.4210 0.6630 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.0890 0.2490 7.2010 0.3590 ;
        RECT 7.1000 0.3590 7.1500 0.5270 ;
        RECT 6.8750 0.5270 7.1500 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5290 0.7050 2.6850 0.7310 ;
        RECT 2.5290 0.7310 2.9890 0.7810 ;
        RECT 2.6350 0.5970 2.6850 0.7050 ;
        RECT 2.5290 0.7810 2.6850 0.8150 ;
        RECT 2.9390 0.7810 2.9890 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 5.5830 0.9420 7.2010 1.0020 ;
        RECT 7.0910 0.6900 7.2010 0.9420 ;
        RECT 6.9670 0.6270 7.0170 0.9420 ;
    END
  END VDDG
  OBS
    LAYER PO ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 2.9490 0.8390 2.9790 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 1.7330 0.7300 1.7630 1.6060 ;
      RECT 3.7090 0.0660 3.7390 0.6910 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 1.2770 0.8400 1.3070 1.6060 ;
      RECT 3.7090 0.9390 3.7390 1.6060 ;
      RECT 3.4050 0.0660 3.4350 0.6370 ;
      RECT 1.2770 0.0660 1.3070 0.6370 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 2.9490 0.0660 2.9790 0.6910 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 2.6450 0.8920 2.6750 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 3.4050 0.8390 3.4350 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 1.7330 0.0680 1.7630 0.6180 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 2.6450 0.0660 2.6750 0.6910 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 4.9250 0.0670 4.9550 1.6050 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
    LAYER NWELL ;
      RECT 5.2800 0.4910 7.2910 1.0830 ;
      RECT -0.1150 1.5430 8.0260 1.7730 ;
      RECT -0.1150 0.6790 4.8180 1.5430 ;
      RECT 7.7510 0.6790 8.0260 1.5430 ;
    LAYER M1 ;
      RECT 4.1390 0.6320 4.5090 0.6820 ;
      RECT 4.4590 0.5970 4.5090 0.6320 ;
      RECT 3.8360 0.4500 3.8860 1.1790 ;
      RECT 3.4720 1.1790 3.9930 1.2290 ;
      RECT 4.2650 0.4500 4.3150 0.6320 ;
      RECT 3.4710 0.4000 4.3150 0.4500 ;
      RECT 3.4710 0.4500 3.5210 0.5630 ;
      RECT 3.4710 0.2970 3.5210 0.4000 ;
      RECT 3.4720 1.2290 3.5220 1.3530 ;
      RECT 4.8990 1.1990 6.1970 1.2490 ;
      RECT 0.4310 1.0830 1.2410 1.1330 ;
      RECT 1.1910 1.1330 1.2410 1.3540 ;
      RECT 1.1910 0.8630 1.2410 1.0830 ;
      RECT 1.1910 0.8130 1.2810 0.8630 ;
      RECT 1.2310 0.4620 1.2810 0.8130 ;
      RECT 1.1750 0.4120 1.2810 0.4620 ;
      RECT 0.4310 0.8690 0.4810 1.0830 ;
      RECT 0.4310 0.8190 0.5210 0.8690 ;
      RECT 0.4310 0.4250 0.5210 0.4750 ;
      RECT 0.4310 0.3620 0.4810 0.4250 ;
      RECT 0.4710 0.4750 0.5210 0.8190 ;
      RECT 3.3190 0.8670 3.4610 0.9170 ;
      RECT 3.3190 0.6630 3.3690 0.8670 ;
      RECT 3.3190 0.6130 3.7650 0.6630 ;
      RECT 3.0190 0.1780 3.6130 0.2280 ;
      RECT 3.0190 0.2280 3.0690 0.2840 ;
      RECT 2.3780 0.2840 3.0690 0.3340 ;
      RECT 1.7230 0.5240 1.7730 0.6130 ;
      RECT 1.9580 0.4550 2.0080 0.6130 ;
      RECT 1.7230 0.6130 2.0080 0.6630 ;
      RECT 2.3780 0.3340 2.4280 0.4050 ;
      RECT 1.9580 0.4050 2.4280 0.4550 ;
      RECT 3.6300 0.9670 3.7650 1.0170 ;
      RECT 3.6300 0.9160 3.6800 0.9670 ;
      RECT 3.5310 0.8660 3.6800 0.9160 ;
      RECT 2.5430 0.4840 3.1040 0.5070 ;
      RECT 2.5430 0.5070 3.1050 0.5340 ;
      RECT 3.0550 0.5340 3.1050 1.0200 ;
      RECT 2.5590 1.0200 3.1050 1.0700 ;
      RECT 2.2950 0.7880 2.3450 1.1200 ;
      RECT 1.5490 0.7380 2.3470 0.7880 ;
      RECT 2.1030 0.5050 2.1530 0.7380 ;
      RECT 2.5590 1.0700 2.6090 1.1200 ;
      RECT 1.9350 1.1200 2.6090 1.1700 ;
      RECT 4.5590 0.6130 4.9810 0.6630 ;
      RECT 4.0030 0.5670 4.0530 0.7590 ;
      RECT 4.2310 0.8090 4.2810 1.3010 ;
      RECT 4.0020 0.5170 4.1450 0.5670 ;
      RECT 4.5590 0.6630 4.6090 0.7590 ;
      RECT 4.0020 0.7590 4.6090 0.8090 ;
      RECT 0.5830 0.6130 1.0290 0.6630 ;
      RECT 0.5830 0.6630 0.6330 1.0040 ;
      RECT 0.5830 0.4130 0.6330 0.6130 ;
      RECT 0.7940 0.0940 1.4910 0.1440 ;
      RECT 5.8870 0.8200 6.4350 0.8700 ;
      RECT 1.3430 0.8540 2.0930 0.9040 ;
      RECT 1.3430 0.4840 1.3930 0.8540 ;
      RECT 1.3430 0.9040 1.3930 1.0990 ;
      RECT 1.3430 0.4340 1.5610 0.4840 ;
      RECT 1.3430 1.0990 1.5610 1.1490 ;
      RECT 1.3430 0.4080 1.3930 0.4340 ;
      RECT 1.3430 1.1490 1.3930 1.3370 ;
      RECT 6.1910 0.7090 6.7290 0.7590 ;
      RECT 1.4030 1.4240 1.7890 1.4740 ;
      RECT 6.8150 0.6770 6.8650 0.7680 ;
      RECT 6.7750 0.4270 6.8650 0.4620 ;
      RECT 6.8150 0.1260 6.8650 0.4270 ;
      RECT 6.7750 0.6270 6.8650 0.6770 ;
      RECT 6.7750 0.5120 6.8250 0.6270 ;
      RECT 6.5710 0.4770 6.8250 0.5120 ;
      RECT 6.5710 0.4620 6.8650 0.4770 ;
      RECT 6.1910 0.1320 6.4250 0.1820 ;
      RECT 5.4470 1.0620 5.8960 1.1120 ;
      RECT 5.4470 0.6770 5.4970 1.0620 ;
      RECT 5.4070 0.6270 5.4970 0.6770 ;
      RECT 5.4070 0.4770 5.4570 0.6270 ;
      RECT 5.4070 0.4270 5.4970 0.4770 ;
      RECT 5.4470 0.1260 5.4970 0.4270 ;
      RECT 1.0990 1.5240 1.9410 1.5740 ;
      RECT 5.5070 0.5270 6.1050 0.5770 ;
      RECT 5.7510 0.5770 5.8010 0.8840 ;
      RECT 5.7510 0.1260 5.8010 0.5270 ;
      RECT 6.0550 0.5770 6.1050 0.7700 ;
      RECT 6.0550 0.3480 6.1050 0.5270 ;
      RECT 3.8350 0.0880 4.0690 0.1380 ;
      RECT 6.4190 1.0620 6.9570 1.1120 ;
      RECT 5.8870 0.2480 6.7290 0.2980 ;
      RECT 3.0730 1.5200 5.8930 1.5700 ;
      RECT 2.3150 1.5200 3.0050 1.5700 ;
      RECT 2.7700 0.6130 3.0050 0.6630 ;
      RECT 2.4070 0.9200 2.8370 0.9700 ;
      RECT 2.7870 0.8310 2.8370 0.9200 ;
      RECT 2.4070 0.9700 2.4570 1.0340 ;
      RECT 2.4070 0.5050 2.4570 0.9200 ;
      RECT 2.1630 1.4200 3.4690 1.4700 ;
      RECT 1.0390 0.7130 1.1650 0.7630 ;
      RECT 1.0390 0.7630 1.0890 1.0330 ;
      RECT 1.1150 0.5630 1.1650 0.7130 ;
      RECT 1.0230 0.5130 1.1650 0.5630 ;
      RECT 2.6950 0.3840 3.3690 0.4340 ;
      RECT 3.3190 0.4340 3.3690 0.5630 ;
      RECT 3.3190 0.2970 3.3690 0.3840 ;
      RECT 3.1670 0.4340 3.2170 0.9670 ;
      RECT 3.1670 0.9670 3.3850 1.0170 ;
      RECT 3.1670 1.0170 3.2170 1.1200 ;
      RECT 3.1670 1.1700 3.2170 1.2700 ;
      RECT 2.6950 1.1200 3.2170 1.1700 ;
      RECT 1.7030 0.9680 2.2150 1.0180 ;
      RECT 2.1620 0.9080 2.2120 0.9680 ;
      RECT 2.1620 0.8580 2.2450 0.9080 ;
  END
END RDFFSRX1_LVT

MACRO RDFFSRX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.208 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 8.2080 1.7020 ;
        RECT 0.2790 1.1310 0.3290 1.6420 ;
        RECT 0.8870 1.2940 0.9370 1.6420 ;
        RECT 1.9910 1.2700 2.0410 1.6420 ;
        RECT 6.2470 1.4540 6.2970 1.6420 ;
        RECT 0.7150 1.2440 0.9370 1.2940 ;
        RECT 1.7830 1.2200 2.9290 1.2700 ;
        RECT 3.6230 1.4040 6.2970 1.4540 ;
        RECT 3.6230 1.2790 3.6730 1.4040 ;
        RECT 4.9910 1.0530 5.0410 1.4040 ;
        RECT 4.6870 0.9610 4.7370 1.4040 ;
        RECT 4.3830 0.9130 4.4330 1.4040 ;
        RECT 4.0790 0.9530 4.1290 1.4040 ;
    END
  END VDD

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6430 1.4650 0.8150 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 8.2080 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.2570 ;
        RECT 4.9910 0.0300 5.0410 0.2210 ;
        RECT 6.8150 0.0300 6.8650 0.1980 ;
        RECT 4.3830 0.0300 4.4330 0.4090 ;
        RECT 4.6870 0.0300 4.7370 0.3200 ;
        RECT 7.2710 0.0300 7.3210 0.4260 ;
        RECT 5.9030 0.0300 5.9530 0.4260 ;
        RECT 4.2550 0.0300 4.3050 0.2830 ;
        RECT 0.2790 0.2570 2.0010 0.3070 ;
        RECT 3.6070 0.2830 4.3050 0.3330 ;
        RECT 0.7350 0.3070 0.7850 0.5570 ;
        RECT 0.8870 0.3070 0.9370 0.5570 ;
        RECT 0.2790 0.3070 0.3290 0.4050 ;
        RECT 1.9510 0.2340 2.0010 0.2570 ;
        RECT 1.9510 0.1840 2.9290 0.2340 ;
        RECT 2.2550 0.2340 2.3050 0.3490 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.4210 0.6630 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2650 0.4010 5.3770 0.4020 ;
        RECT 4.5350 0.4020 5.3870 0.4520 ;
        RECT 4.5350 0.1490 4.5850 0.4020 ;
        RECT 5.2650 0.4520 5.3870 0.5120 ;
        RECT 5.3370 0.5120 5.3870 0.8330 ;
        RECT 4.5350 0.8330 5.3870 0.8830 ;
        RECT 4.5350 0.8830 4.5850 1.3190 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8390 0.1490 4.8890 0.2710 ;
        RECT 4.8390 0.2710 5.5370 0.3210 ;
        RECT 5.4170 0.3210 5.5370 0.3600 ;
        RECT 5.4170 0.2500 5.5370 0.2710 ;
        RECT 5.4870 0.3600 5.5370 0.9330 ;
        RECT 5.4170 0.2490 5.5290 0.2500 ;
        RECT 4.8390 0.9330 5.5370 0.9830 ;
        RECT 4.8390 0.9830 4.8890 1.3270 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.3930 0.2490 7.5050 0.3590 ;
        RECT 7.4040 0.3590 7.4540 0.5270 ;
        RECT 7.1790 0.5270 7.4540 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5290 0.7050 2.6850 0.7310 ;
        RECT 2.5290 0.7310 2.9890 0.7810 ;
        RECT 2.6350 0.5970 2.6850 0.7050 ;
        RECT 2.5290 0.7810 2.6850 0.8150 ;
        RECT 2.9390 0.7810 2.9890 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 5.8870 0.9420 7.5050 1.0020 ;
        RECT 7.3950 0.6900 7.5050 0.9420 ;
        RECT 7.2710 0.6270 7.3210 0.9420 ;
    END
  END VDDG
  OBS
    LAYER PO ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 2.9490 0.8390 2.9790 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 1.7330 0.7300 1.7630 1.6060 ;
      RECT 3.7090 0.0660 3.7390 0.6910 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 1.2770 0.8400 1.3070 1.6060 ;
      RECT 3.7090 0.9390 3.7390 1.6060 ;
      RECT 3.4050 0.0660 3.4350 0.6370 ;
      RECT 1.2770 0.0660 1.3070 0.6370 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 2.9490 0.0660 2.9790 0.6910 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 2.6450 0.8920 2.6750 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
      RECT 3.4050 0.8390 3.4350 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 1.7330 0.0680 1.7630 0.6180 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 2.6450 0.0660 2.6750 0.6910 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 5.2290 0.0670 5.2590 1.6050 ;
    LAYER NWELL ;
      RECT 5.5840 0.4910 7.5950 1.0830 ;
      RECT -0.1150 1.5430 8.3300 1.7730 ;
      RECT -0.1150 0.6790 5.1220 1.5430 ;
      RECT 8.0550 0.6790 8.3300 1.5430 ;
    LAYER M1 ;
      RECT 4.1390 0.6320 4.6770 0.6820 ;
      RECT 3.4710 0.4500 3.5210 0.5630 ;
      RECT 3.4710 0.2970 3.5210 0.4000 ;
      RECT 3.4720 1.2290 3.5220 1.3530 ;
      RECT 3.8360 0.4500 3.8860 1.1790 ;
      RECT 3.4720 1.1790 3.9930 1.2290 ;
      RECT 3.4710 0.4000 4.3150 0.4500 ;
      RECT 4.2650 0.4500 4.3150 0.6320 ;
      RECT 1.0390 0.7130 1.1650 0.7630 ;
      RECT 1.0390 0.7630 1.0890 1.0330 ;
      RECT 1.1150 0.5630 1.1650 0.7130 ;
      RECT 1.0230 0.5130 1.1650 0.5630 ;
      RECT 2.6950 0.3840 3.3690 0.4340 ;
      RECT 3.3190 0.4340 3.3690 0.5630 ;
      RECT 3.3190 0.2970 3.3690 0.3840 ;
      RECT 3.1670 0.4340 3.2170 0.9670 ;
      RECT 3.1670 0.9670 3.3850 1.0170 ;
      RECT 3.1670 1.0170 3.2170 1.1200 ;
      RECT 3.1670 1.1700 3.2170 1.2700 ;
      RECT 2.6950 1.1200 3.2170 1.1700 ;
      RECT 1.7030 0.9680 2.2150 1.0180 ;
      RECT 2.1620 0.9080 2.2120 0.9680 ;
      RECT 2.1620 0.8580 2.2450 0.9080 ;
      RECT 4.7270 0.6130 5.2850 0.6630 ;
      RECT 4.0030 0.7820 4.0530 0.8090 ;
      RECT 4.0030 0.5670 4.0530 0.7320 ;
      RECT 4.2310 0.7820 4.2810 1.3010 ;
      RECT 4.0020 0.5170 4.1450 0.5670 ;
      RECT 4.7270 0.6630 4.7770 0.7320 ;
      RECT 4.0020 0.7320 4.7770 0.7820 ;
      RECT 3.3190 0.8670 3.4610 0.9170 ;
      RECT 3.3190 0.6630 3.3690 0.8670 ;
      RECT 3.3190 0.6130 3.7650 0.6630 ;
      RECT 3.0190 0.1780 3.6130 0.2280 ;
      RECT 3.0190 0.2280 3.0690 0.2840 ;
      RECT 2.3780 0.2840 3.0690 0.3340 ;
      RECT 1.7230 0.5240 1.7730 0.6130 ;
      RECT 1.9580 0.4550 2.0080 0.6130 ;
      RECT 1.7230 0.6130 2.0080 0.6630 ;
      RECT 2.3780 0.3340 2.4280 0.4050 ;
      RECT 1.9580 0.4050 2.4280 0.4550 ;
      RECT 2.4070 0.9200 2.8370 0.9700 ;
      RECT 2.7870 0.8310 2.8370 0.9200 ;
      RECT 2.4070 0.9700 2.4570 1.0340 ;
      RECT 2.4070 0.5050 2.4570 0.9200 ;
      RECT 2.1630 1.4200 3.4690 1.4700 ;
      RECT 1.1910 0.8130 1.2810 0.8630 ;
      RECT 1.1910 0.8630 1.2410 1.0830 ;
      RECT 1.2310 0.4620 1.2810 0.8130 ;
      RECT 0.4310 1.0830 1.2410 1.1330 ;
      RECT 1.1750 0.4120 1.2810 0.4620 ;
      RECT 1.1910 1.1330 1.2410 1.3540 ;
      RECT 0.4310 0.8690 0.4810 1.0830 ;
      RECT 0.4310 0.8190 0.5210 0.8690 ;
      RECT 0.4310 0.4250 0.5210 0.4750 ;
      RECT 0.4310 0.3620 0.4810 0.4250 ;
      RECT 0.4710 0.4750 0.5210 0.8190 ;
      RECT 5.2030 1.1990 6.5010 1.2490 ;
      RECT 3.6300 0.9670 3.7650 1.0170 ;
      RECT 3.6300 0.9160 3.6800 0.9670 ;
      RECT 3.5310 0.8660 3.6800 0.9160 ;
      RECT 2.5430 0.4840 3.1040 0.5070 ;
      RECT 2.5430 0.5070 3.1050 0.5340 ;
      RECT 3.0550 0.5340 3.1050 1.0200 ;
      RECT 2.5590 1.0200 3.1050 1.0700 ;
      RECT 2.2950 0.7880 2.3450 1.1200 ;
      RECT 1.5490 0.7380 2.3470 0.7880 ;
      RECT 2.1030 0.5050 2.1530 0.7380 ;
      RECT 2.5590 1.0700 2.6090 1.1200 ;
      RECT 1.9350 1.1200 2.6090 1.1700 ;
      RECT 0.5830 0.6130 1.0290 0.6630 ;
      RECT 0.5830 0.6630 0.6330 1.0040 ;
      RECT 0.5830 0.4130 0.6330 0.6130 ;
      RECT 0.7940 0.0940 1.4910 0.1440 ;
      RECT 6.1910 0.8200 6.7390 0.8700 ;
      RECT 1.3430 0.8540 2.0930 0.9040 ;
      RECT 1.3430 0.4840 1.3930 0.8540 ;
      RECT 1.3430 0.9040 1.3930 1.0990 ;
      RECT 1.3430 0.4340 1.5610 0.4840 ;
      RECT 1.3430 1.0990 1.5610 1.1490 ;
      RECT 1.3430 0.4080 1.3930 0.4340 ;
      RECT 1.3430 1.1490 1.3930 1.3370 ;
      RECT 6.4950 0.7090 7.0330 0.7590 ;
      RECT 1.4030 1.4240 1.7890 1.4740 ;
      RECT 7.1190 0.6770 7.1690 0.7680 ;
      RECT 7.0790 0.4270 7.1690 0.4620 ;
      RECT 7.1190 0.1260 7.1690 0.4270 ;
      RECT 7.0790 0.6270 7.1690 0.6770 ;
      RECT 7.0790 0.5120 7.1290 0.6270 ;
      RECT 6.8750 0.4770 7.1290 0.5120 ;
      RECT 6.8750 0.4620 7.1690 0.4770 ;
      RECT 6.4950 0.1320 6.7290 0.1820 ;
      RECT 5.7510 1.0620 6.2000 1.1120 ;
      RECT 5.7510 0.6770 5.8010 1.0620 ;
      RECT 5.7110 0.6270 5.8010 0.6770 ;
      RECT 5.7110 0.4770 5.7610 0.6270 ;
      RECT 5.7110 0.4270 5.8010 0.4770 ;
      RECT 5.7510 0.1260 5.8010 0.4270 ;
      RECT 1.0990 1.5240 1.9410 1.5740 ;
      RECT 5.8110 0.5270 6.4090 0.5770 ;
      RECT 6.0550 0.5770 6.1050 0.8840 ;
      RECT 6.0550 0.1260 6.1050 0.5270 ;
      RECT 6.3590 0.5770 6.4090 0.7700 ;
      RECT 6.3590 0.3480 6.4090 0.5270 ;
      RECT 3.8350 0.0880 4.0690 0.1380 ;
      RECT 6.7230 1.0620 7.2610 1.1120 ;
      RECT 6.1910 0.2480 7.0330 0.2980 ;
      RECT 3.0730 1.5200 6.1970 1.5700 ;
      RECT 2.3150 1.5200 3.0050 1.5700 ;
      RECT 2.7700 0.6130 3.0050 0.6630 ;
  END
END RDFFSRX2_LVT

MACRO RDFFX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.36 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 6.1910 0.9420 7.6580 1.0020 ;
        RECT 7.5480 0.6900 7.6580 0.9420 ;
    END
  END VDDG

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 8.3600 0.0300 ;
        RECT 0.5830 0.0300 0.6330 0.3070 ;
        RECT 7.2710 0.0300 7.3210 0.3120 ;
        RECT 0.4310 0.0300 0.4810 0.5570 ;
        RECT 5.1430 0.0300 5.1930 0.2410 ;
        RECT 6.9670 0.0300 7.0170 0.2020 ;
        RECT 6.2070 0.0300 6.2570 0.2060 ;
        RECT 4.8790 0.0300 4.9290 0.2830 ;
        RECT 0.5830 0.3070 2.1530 0.3570 ;
        RECT 2.9990 0.2830 4.9300 0.3330 ;
        RECT 1.4950 0.3570 1.5450 0.5580 ;
        RECT 1.6470 0.3570 1.6970 0.5580 ;
        RECT 2.1030 0.3570 2.1530 0.5770 ;
        RECT 4.8390 0.3330 4.8890 0.4430 ;
    END
  END VSS

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 1.4650 0.4220 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2950 0.9690 5.8290 1.0190 ;
        RECT 5.7790 0.3510 5.8290 0.9690 ;
        RECT 5.2950 1.0190 5.5270 1.1290 ;
        RECT 5.2790 0.3010 5.8290 0.3510 ;
        RECT 5.2950 1.1290 5.3450 1.3270 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.9910 0.1570 5.0410 0.4010 ;
        RECT 4.9910 0.4010 5.6910 0.4510 ;
        RECT 5.5690 0.4510 5.6910 0.5380 ;
        RECT 5.6410 0.5380 5.6910 0.8590 ;
        RECT 4.9910 0.8590 5.6910 0.9090 ;
        RECT 4.9910 0.9090 5.0410 1.2320 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 8.3600 1.7020 ;
        RECT 0.5430 1.3400 0.5930 1.6420 ;
        RECT 3.2070 1.3400 3.2570 1.6420 ;
        RECT 0.4130 1.2900 5.1940 1.3400 ;
        RECT 3.0150 0.9730 3.0650 1.2900 ;
        RECT 5.1430 0.9590 5.1930 1.2900 ;
    END
  END VDD

  PIN RETN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.5130 1.4080 6.8980 1.4580 ;
        RECT 6.7850 1.3130 6.8980 1.4080 ;
    END
    ANTENNAGATEAREA 0.084 ;
  END RETN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0970 0.9670 1.1810 1.0170 ;
        RECT 0.0970 1.0170 0.2080 1.1190 ;
    END
    ANTENNAGATEAREA 0.018 ;
  END D
  OBS
    LAYER PO ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 3.5570 0.9590 3.5870 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 5.5330 0.0670 5.5630 1.6050 ;
      RECT 1.7330 0.9390 1.7630 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 1.7330 0.0660 1.7630 0.6370 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 0.9730 0.0660 1.0030 0.6910 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 2.1890 0.9390 2.2190 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 3.5570 0.0660 3.5870 0.6910 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 4.0130 0.0660 4.0430 0.7910 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 2.6450 0.0660 2.6750 0.6910 ;
      RECT 2.1890 0.0660 2.2190 0.6370 ;
      RECT 0.9730 0.8390 1.0030 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 4.0130 0.9390 4.0430 1.6060 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 2.6450 0.8390 2.6750 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 3.7090 0.0660 3.7390 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
    LAYER NWELL ;
      RECT -0.1160 1.5430 8.4690 1.7730 ;
      RECT -0.1160 0.6790 5.4270 1.5430 ;
      RECT 8.1950 0.6790 8.4690 1.5430 ;
      RECT 5.8890 0.4910 7.7350 1.0830 ;
    LAYER M1 ;
      RECT 7.2620 0.4120 7.3120 0.4620 ;
      RECT 7.2620 0.4620 7.4130 0.5120 ;
      RECT 7.2620 0.5120 7.3120 0.5890 ;
      RECT 7.1190 0.5890 7.3120 0.6390 ;
      RECT 7.1190 0.3620 7.3120 0.4120 ;
      RECT 7.1190 0.1260 7.1690 0.3620 ;
      RECT 7.1190 0.6390 7.1690 0.7820 ;
      RECT 1.9110 0.8670 2.1930 0.9170 ;
      RECT 2.1430 0.9170 2.1930 1.1270 ;
      RECT 1.1910 1.1270 2.1930 1.1770 ;
      RECT 1.1910 1.1770 1.2410 1.2400 ;
      RECT 1.2410 0.9170 1.2910 1.0660 ;
      RECT 1.1910 0.4130 1.2410 0.8670 ;
      RECT 1.9110 0.6070 1.9610 0.8670 ;
      RECT 1.9110 0.5570 2.0010 0.6070 ;
      RECT 1.9510 0.4130 2.0010 0.5570 ;
      RECT 1.1910 1.0670 1.2910 1.1270 ;
      RECT 1.2310 1.0660 1.2910 1.0670 ;
      RECT 1.1910 0.8670 1.4850 0.9170 ;
      RECT 2.8230 0.7670 2.9530 0.8170 ;
      RECT 2.9030 0.5630 2.9530 0.7670 ;
      RECT 2.8630 0.5130 2.9530 0.5630 ;
      RECT 2.7110 1.1900 2.9130 1.2400 ;
      RECT 2.7110 0.9740 2.7610 1.1900 ;
      RECT 2.8630 1.0240 2.9130 1.1900 ;
      RECT 2.8230 0.9740 2.9130 1.0240 ;
      RECT 2.8230 0.8170 2.8730 0.9740 ;
      RECT 2.8630 0.3270 2.9130 0.5130 ;
      RECT 2.7110 0.2770 2.9130 0.3270 ;
      RECT 2.7110 0.3270 2.7610 0.5560 ;
      RECT 0.6430 1.5240 2.8530 1.5740 ;
      RECT 0.7950 0.0940 2.5490 0.1440 ;
      RECT 3.1270 0.7670 3.3690 0.8170 ;
      RECT 3.3190 0.8170 3.3690 1.2400 ;
      RECT 3.1270 0.4530 3.1770 0.7670 ;
      RECT 3.0030 0.4030 3.3700 0.4530 ;
      RECT 3.3190 0.4530 3.3690 0.5770 ;
      RECT 3.0030 0.4530 3.0530 0.8670 ;
      RECT 2.9230 0.8670 3.0530 0.9170 ;
      RECT 3.4310 0.5130 4.2970 0.5630 ;
      RECT 3.4310 0.5630 3.4810 0.6270 ;
      RECT 3.2270 0.6270 3.4810 0.6770 ;
      RECT 3.4310 0.6770 3.4810 1.0670 ;
      RECT 3.4310 1.0670 4.2970 1.1170 ;
      RECT 3.5310 0.6130 4.4330 0.6630 ;
      RECT 4.3830 0.3830 4.4330 0.6130 ;
      RECT 3.7350 0.6630 3.7850 0.9670 ;
      RECT 3.7350 0.9670 4.4330 1.0170 ;
      RECT 4.3830 1.0170 4.4330 1.2400 ;
      RECT 6.8150 0.4620 7.1090 0.5120 ;
      RECT 6.8150 0.1820 6.8650 0.4620 ;
      RECT 6.8150 0.5120 6.8650 0.6350 ;
      RECT 6.4950 0.1320 6.8650 0.1820 ;
      RECT 6.4950 0.6350 6.8650 0.6850 ;
      RECT 6.3590 0.4940 6.7130 0.5440 ;
      RECT 6.6630 0.3480 6.7130 0.4940 ;
      RECT 6.3590 0.5440 6.4090 0.7820 ;
      RECT 4.1390 0.7590 5.5890 0.8090 ;
      RECT 5.0670 0.6420 5.1170 0.7590 ;
      RECT 4.6870 0.8090 4.7370 1.2400 ;
      RECT 4.4950 0.5630 4.5450 0.7590 ;
      RECT 4.4950 0.5130 4.7370 0.5630 ;
      RECT 4.6870 0.3830 4.7370 0.5130 ;
      RECT 3.6830 1.5280 7.7190 1.5780 ;
      RECT 3.8350 0.7130 4.0690 0.7630 ;
      RECT 1.4790 0.9670 2.0930 1.0170 ;
      RECT 1.3430 0.4070 1.3930 0.6190 ;
      RECT 1.6470 0.6690 1.6970 0.9670 ;
      RECT 1.3430 0.6190 1.6970 0.6690 ;
      RECT 7.4230 0.5620 7.7170 0.6120 ;
      RECT 7.5580 0.4120 7.6080 0.5620 ;
      RECT 7.4230 0.3620 7.6080 0.4120 ;
      RECT 7.4230 0.6120 7.4730 0.8320 ;
      RECT 6.2590 0.8320 7.4730 0.8820 ;
      RECT 7.4230 0.1260 7.4730 0.3620 ;
      RECT 6.2590 0.4200 6.3090 0.8320 ;
      RECT 6.2590 0.3700 6.4270 0.4200 ;
      RECT 2.4670 0.8670 2.7210 0.9170 ;
      RECT 0.2790 0.6130 0.7250 0.6630 ;
      RECT 0.6090 0.4630 0.6590 0.6130 ;
      RECT 0.6090 0.4130 1.0130 0.4630 ;
      RECT 0.9630 0.4630 1.0130 0.6800 ;
      RECT 0.2790 0.6630 0.3290 0.9120 ;
      RECT 0.2790 0.4130 0.3290 0.6130 ;
      RECT 0.7190 0.5130 0.8610 0.5630 ;
      RECT 0.8110 0.5630 0.8610 0.7130 ;
      RECT 0.7350 0.7130 0.8610 0.7630 ;
      RECT 0.7350 0.7630 0.7850 0.8670 ;
      RECT 0.7350 0.8670 1.0290 0.9170 ;
      RECT 2.0110 0.6670 2.3970 0.7170 ;
      RECT 5.5070 1.2000 6.6530 1.2500 ;
      RECT 2.6190 0.6130 2.8530 0.6630 ;
      RECT 4.9670 0.5010 5.2690 0.5510 ;
      RECT 5.2190 0.5510 5.2690 0.6790 ;
      RECT 4.9670 0.5510 5.0170 0.6130 ;
      RECT 4.5950 0.6130 5.0170 0.6630 ;
      RECT 6.0550 1.0620 6.5010 1.1120 ;
      RECT 6.0550 0.1260 6.1050 1.0620 ;
      RECT 2.5990 0.0920 4.6780 0.1420 ;
      RECT 2.5990 0.1420 2.6490 0.1940 ;
      RECT 2.5590 0.1940 2.6490 0.2440 ;
      RECT 2.5590 0.2440 2.6090 0.5130 ;
      RECT 2.4070 0.5130 2.6090 0.5630 ;
      RECT 2.4070 0.2770 2.4570 0.5130 ;
      RECT 2.4470 0.5630 2.4970 0.7670 ;
      RECT 2.3670 0.7670 2.4970 0.8170 ;
      RECT 2.3670 0.8170 2.4170 0.9670 ;
      RECT 2.3670 0.9670 2.4570 1.0170 ;
      RECT 2.4070 1.0170 2.4570 1.1900 ;
      RECT 2.4070 1.1900 2.6090 1.2400 ;
      RECT 2.5590 0.9740 2.6090 1.1900 ;
  END
END RDFFX1_LVT

MACRO RDFFX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.664 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 6.4950 0.9420 7.9620 1.0020 ;
        RECT 7.8520 0.6900 7.9620 0.9420 ;
    END
  END VDDG

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 8.6640 0.0300 ;
        RECT 0.5830 0.0300 0.6330 0.3070 ;
        RECT 7.5750 0.0300 7.6250 0.3120 ;
        RECT 6.5110 0.0300 6.5610 0.2060 ;
        RECT 0.4310 0.0300 0.4810 0.5570 ;
        RECT 5.5990 0.0300 5.6490 0.2210 ;
        RECT 5.2950 0.0300 5.3450 0.3200 ;
        RECT 7.2710 0.0300 7.3210 0.2020 ;
        RECT 4.9910 0.0300 5.0410 0.2830 ;
        RECT 0.5830 0.3070 2.1530 0.3570 ;
        RECT 2.9990 0.2830 5.0410 0.3330 ;
        RECT 2.1030 0.3570 2.1530 0.5770 ;
        RECT 1.4950 0.3570 1.5450 0.5580 ;
        RECT 1.6470 0.3570 1.6970 0.5580 ;
        RECT 4.8390 0.3330 4.8890 0.4430 ;
        RECT 4.9910 0.3330 5.0410 0.4090 ;
    END
  END VSS

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 1.4650 0.4220 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 8.6640 1.7020 ;
        RECT 0.5430 1.3400 0.5930 1.6420 ;
        RECT 3.2070 1.3400 3.2570 1.6420 ;
        RECT 0.4130 1.2900 5.6490 1.3400 ;
        RECT 5.5990 1.0530 5.6490 1.2900 ;
        RECT 5.2950 0.9610 5.3450 1.2900 ;
        RECT 3.0150 0.9730 3.0650 1.2900 ;
        RECT 4.9910 0.9130 5.0410 1.2900 ;
    END
  END VDD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4470 0.1490 5.4970 0.2710 ;
        RECT 5.4470 0.2710 6.1450 0.3210 ;
        RECT 6.0250 0.3210 6.1450 0.3590 ;
        RECT 6.0250 0.2500 6.1450 0.2710 ;
        RECT 6.0950 0.3590 6.1450 0.9330 ;
        RECT 6.0250 0.2490 6.1370 0.2500 ;
        RECT 5.4470 0.9330 6.1450 0.9830 ;
        RECT 5.4470 0.9830 5.4970 1.2240 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8730 0.4010 5.9850 0.4020 ;
        RECT 5.1430 0.4020 5.9950 0.4520 ;
        RECT 5.1430 0.1490 5.1930 0.4020 ;
        RECT 5.8730 0.4520 5.9950 0.5120 ;
        RECT 5.9450 0.5120 5.9950 0.8330 ;
        RECT 5.1430 0.8330 5.9950 0.8830 ;
        RECT 5.1430 0.8830 5.1930 1.2240 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN RETN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.5130 1.4080 7.2020 1.4580 ;
        RECT 7.0890 1.3130 7.2020 1.4080 ;
    END
    ANTENNAGATEAREA 0.084 ;
  END RETN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0970 0.9670 1.1810 1.0170 ;
        RECT 0.0970 1.0170 0.2080 1.1190 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D
  OBS
    LAYER PO ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 3.7090 0.0660 3.7390 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 3.5570 0.9590 3.5870 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 5.8370 0.0670 5.8670 1.6050 ;
      RECT 1.7330 0.9390 1.7630 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 1.7330 0.0660 1.7630 0.6370 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 0.9730 0.0660 1.0030 0.6910 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 2.1890 0.9390 2.2190 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 3.5570 0.0660 3.5870 0.6910 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 4.0130 0.0660 4.0430 0.7910 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 2.6450 0.0660 2.6750 0.6910 ;
      RECT 2.1890 0.0660 2.2190 0.6370 ;
      RECT 0.9730 0.8390 1.0030 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 4.0130 0.9390 4.0430 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 2.6450 0.8390 2.6750 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
    LAYER NWELL ;
      RECT -0.1160 1.5430 8.7740 1.7730 ;
      RECT -0.1160 0.6790 5.7310 1.5430 ;
      RECT 8.4990 0.6790 8.7740 1.5430 ;
      RECT 6.1930 0.4910 8.0390 1.0830 ;
    LAYER M1 ;
      RECT 2.5990 0.0920 4.6780 0.1420 ;
      RECT 2.4070 0.2770 2.4570 0.5130 ;
      RECT 2.4070 0.5130 2.6090 0.5630 ;
      RECT 2.5590 0.2440 2.6090 0.5130 ;
      RECT 2.4470 0.5630 2.4970 0.7670 ;
      RECT 2.5590 0.1940 2.6490 0.2440 ;
      RECT 2.3670 0.7670 2.4970 0.8170 ;
      RECT 2.5990 0.1420 2.6490 0.1940 ;
      RECT 2.3670 0.8170 2.4170 0.9670 ;
      RECT 2.3670 0.9670 2.4570 1.0170 ;
      RECT 2.4070 1.0170 2.4570 1.1900 ;
      RECT 2.4070 1.1900 2.6090 1.2400 ;
      RECT 2.5590 0.9740 2.6090 1.1900 ;
      RECT 1.9110 0.8670 2.1930 0.9170 ;
      RECT 2.1430 0.9170 2.1930 1.1270 ;
      RECT 1.1910 1.1270 2.1930 1.1770 ;
      RECT 1.1910 1.1770 1.2410 1.2400 ;
      RECT 1.2410 0.9170 1.2910 1.0660 ;
      RECT 1.1910 0.4130 1.2410 0.8670 ;
      RECT 1.9110 0.6070 1.9610 0.8670 ;
      RECT 1.9110 0.5570 2.0010 0.6070 ;
      RECT 1.9510 0.4130 2.0010 0.5570 ;
      RECT 1.1910 1.0670 1.2910 1.1270 ;
      RECT 1.2310 1.0660 1.2910 1.0670 ;
      RECT 1.1910 0.8670 1.4850 0.9170 ;
      RECT 4.1390 0.7130 5.8930 0.7630 ;
      RECT 4.6870 0.7630 4.7370 1.2400 ;
      RECT 4.4950 0.5630 4.5450 0.7130 ;
      RECT 4.4950 0.5130 4.7370 0.5630 ;
      RECT 4.6870 0.3830 4.7370 0.5130 ;
      RECT 5.0670 0.6420 5.1170 0.7130 ;
      RECT 5.2190 0.6420 5.2690 0.7130 ;
      RECT 1.4790 0.9670 2.0930 1.0170 ;
      RECT 1.3430 0.4070 1.3930 0.6190 ;
      RECT 1.6470 0.6690 1.6970 0.9670 ;
      RECT 1.3430 0.6190 1.6970 0.6690 ;
      RECT 2.8630 0.5130 2.9530 0.5630 ;
      RECT 2.9030 0.5630 2.9530 0.7670 ;
      RECT 2.8230 0.7670 2.9530 0.8170 ;
      RECT 2.7110 0.2770 2.9130 0.3270 ;
      RECT 2.7110 0.3270 2.7610 0.5560 ;
      RECT 2.8630 0.3270 2.9130 0.5130 ;
      RECT 2.8230 0.8170 2.8730 0.9740 ;
      RECT 2.8230 0.9740 2.9130 1.0240 ;
      RECT 2.8630 1.0240 2.9130 1.1900 ;
      RECT 2.7110 1.1900 2.9130 1.2400 ;
      RECT 2.7110 0.9740 2.7610 1.1900 ;
      RECT 7.4230 0.5890 7.6160 0.6390 ;
      RECT 7.5660 0.5120 7.6160 0.5890 ;
      RECT 7.5660 0.4620 7.7170 0.5120 ;
      RECT 7.5660 0.4120 7.6160 0.4620 ;
      RECT 7.4230 0.3620 7.6160 0.4120 ;
      RECT 7.4230 0.6390 7.4730 0.7820 ;
      RECT 7.4230 0.1260 7.4730 0.3620 ;
      RECT 2.6190 0.6130 2.8530 0.6630 ;
      RECT 0.6430 1.5240 2.8530 1.5740 ;
      RECT 0.7950 0.0940 2.5490 0.1440 ;
      RECT 3.1270 0.7670 3.3690 0.8170 ;
      RECT 3.3190 0.8170 3.3690 1.2400 ;
      RECT 3.1270 0.4530 3.1770 0.7670 ;
      RECT 3.0030 0.4030 3.3700 0.4530 ;
      RECT 3.3190 0.4530 3.3690 0.5770 ;
      RECT 3.0030 0.4530 3.0530 0.8670 ;
      RECT 2.9230 0.8670 3.0530 0.9170 ;
      RECT 3.4310 0.5130 4.2970 0.5630 ;
      RECT 3.4310 0.5630 3.4810 0.6270 ;
      RECT 3.2270 0.6270 3.4810 0.6770 ;
      RECT 3.4310 0.6770 3.4810 1.0670 ;
      RECT 3.4310 1.0670 4.2970 1.1170 ;
      RECT 3.5310 0.6130 4.4330 0.6630 ;
      RECT 4.3830 0.3830 4.4330 0.6130 ;
      RECT 3.7350 0.6630 3.7850 0.9670 ;
      RECT 3.7350 0.9670 4.4330 1.0170 ;
      RECT 4.3830 1.0170 4.4330 1.2400 ;
      RECT 7.1190 0.4620 7.4130 0.5120 ;
      RECT 7.1190 0.1820 7.1690 0.4620 ;
      RECT 7.1190 0.5120 7.1690 0.6350 ;
      RECT 6.7990 0.1320 7.1690 0.1820 ;
      RECT 6.7990 0.6350 7.1690 0.6850 ;
      RECT 6.6630 0.4940 7.0170 0.5440 ;
      RECT 6.9670 0.3480 7.0170 0.4940 ;
      RECT 6.6630 0.5440 6.7130 0.7820 ;
      RECT 3.6830 1.5280 8.0230 1.5780 ;
      RECT 3.8350 0.7130 4.0690 0.7630 ;
      RECT 7.7270 0.5620 8.0210 0.6120 ;
      RECT 7.8620 0.4120 7.9120 0.5620 ;
      RECT 7.7270 0.3620 7.9120 0.4120 ;
      RECT 7.7270 0.6120 7.7770 0.8320 ;
      RECT 6.5630 0.8320 7.7770 0.8820 ;
      RECT 7.7270 0.1260 7.7770 0.3620 ;
      RECT 6.5630 0.4200 6.6130 0.8320 ;
      RECT 6.5630 0.3700 6.7310 0.4200 ;
      RECT 2.4670 0.8670 2.7210 0.9170 ;
      RECT 0.2790 0.6130 0.7250 0.6630 ;
      RECT 0.6090 0.4630 0.6590 0.6130 ;
      RECT 0.6090 0.4130 1.0130 0.4630 ;
      RECT 0.9630 0.4630 1.0130 0.6800 ;
      RECT 0.2790 0.6630 0.3290 0.9120 ;
      RECT 0.2790 0.4130 0.3290 0.6130 ;
      RECT 0.7190 0.5130 0.8610 0.5630 ;
      RECT 0.8110 0.5630 0.8610 0.7130 ;
      RECT 0.7350 0.7130 0.8610 0.7630 ;
      RECT 0.7350 0.7630 0.7850 0.8670 ;
      RECT 0.7350 0.8670 1.0290 0.9170 ;
      RECT 2.0110 0.6670 2.3970 0.7170 ;
      RECT 5.8110 1.2000 6.9570 1.2500 ;
      RECT 4.9180 0.5200 5.4030 0.5700 ;
      RECT 5.3530 0.5700 5.4030 0.6040 ;
      RECT 4.9180 0.5700 4.9680 0.6130 ;
      RECT 5.3530 0.6040 5.5890 0.6540 ;
      RECT 4.5950 0.6130 4.9680 0.6630 ;
      RECT 6.3590 1.0620 6.8050 1.1120 ;
      RECT 6.3590 0.1260 6.4090 1.0620 ;
  END
END RDFFX2_LVT

MACRO RSDFFARX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.792 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 1.1610 1.0110 1.3160 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6780 0.7250 0.7280 ;
        RECT 0.4010 0.5510 0.5110 0.6780 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 0.0970 1.3180 0.2070 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 8.6230 0.9420 10.0900 1.0020 ;
        RECT 9.9800 0.6900 10.0900 0.9420 ;
    END
  END VDDG

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 10.7920 0.0300 ;
        RECT 2.4070 0.0300 2.4570 0.3070 ;
        RECT 9.7030 0.0300 9.7530 0.3120 ;
        RECT 1.7990 0.0300 1.8490 0.4050 ;
        RECT 9.3990 0.0300 9.4490 0.2020 ;
        RECT 0.4310 0.0300 0.4810 0.4340 ;
        RECT 0.5830 0.0300 0.6330 0.5120 ;
        RECT 8.6390 0.0300 8.6890 0.2060 ;
        RECT 2.2550 0.0300 2.3050 0.5570 ;
        RECT 7.5750 0.0300 7.6250 0.2410 ;
        RECT 1.6470 0.0300 1.6970 0.4050 ;
        RECT 7.3110 0.0300 7.3610 0.2830 ;
        RECT 2.4070 0.3070 4.1290 0.3570 ;
        RECT 4.9750 0.2830 7.3610 0.3330 ;
        RECT 4.0790 0.3570 4.1290 0.5770 ;
        RECT 3.3190 0.3570 3.3690 0.5580 ;
        RECT 3.6230 0.3570 3.6730 0.5580 ;
        RECT 7.2710 0.3330 7.3210 0.4430 ;
    END
  END VSS

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0720 1.4650 2.2460 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.7270 0.9690 8.2610 1.0190 ;
        RECT 7.7270 1.0190 7.9590 1.1290 ;
        RECT 8.2110 0.3510 8.2610 0.9690 ;
        RECT 7.7270 1.1290 7.7770 1.3270 ;
        RECT 7.7110 0.3010 8.2610 0.3510 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.4230 0.1570 7.4730 0.4010 ;
        RECT 7.4230 0.4010 8.1230 0.4510 ;
        RECT 8.0010 0.4510 8.1230 0.5380 ;
        RECT 8.0730 0.5380 8.1230 0.8590 ;
        RECT 7.4230 0.8590 8.1230 0.9090 ;
        RECT 7.4230 0.9090 7.4730 1.2320 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 10.7920 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 1.7990 1.1310 1.8490 1.6420 ;
        RECT 1.6470 1.1310 1.6970 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 5.6390 1.3400 5.6890 1.6420 ;
        RECT 2.3670 1.3400 2.4170 1.6420 ;
        RECT 2.2370 1.2900 7.6250 1.3400 ;
        RECT 7.5750 0.9590 7.6250 1.2900 ;
        RECT 4.9910 0.9730 5.0410 1.2900 ;
    END
  END VDD

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.1130 0.8510 5.2680 0.9670 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END RSTB

  PIN RETN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.9450 1.4080 9.3300 1.4580 ;
        RECT 9.2170 1.3130 9.3300 1.4080 ;
    END
    ANTENNAGATEAREA 0.084 ;
  END RETN
  OBS
    LAYER M1 ;
      RECT 4.3430 0.9670 4.4330 1.0170 ;
      RECT 4.3830 1.0170 4.4330 1.1900 ;
      RECT 4.3830 1.1900 4.5850 1.2400 ;
      RECT 4.5350 0.9740 4.5850 1.1900 ;
      RECT 9.5510 0.5890 9.7440 0.6390 ;
      RECT 9.6940 0.5120 9.7440 0.5890 ;
      RECT 9.6940 0.4620 9.8450 0.5120 ;
      RECT 9.6940 0.4120 9.7440 0.4620 ;
      RECT 9.5510 0.3620 9.7440 0.4120 ;
      RECT 9.5510 0.6390 9.6010 0.7820 ;
      RECT 9.5510 0.1260 9.6010 0.3620 ;
      RECT 8.7910 0.4940 9.1450 0.5440 ;
      RECT 9.0950 0.3480 9.1450 0.4940 ;
      RECT 8.7910 0.5440 8.8410 0.7820 ;
      RECT 9.2470 0.4620 9.5410 0.5120 ;
      RECT 9.2470 0.5120 9.2970 0.6350 ;
      RECT 9.2470 0.1820 9.2970 0.4620 ;
      RECT 8.9270 0.6350 9.2970 0.6850 ;
      RECT 8.9270 0.1320 9.2970 0.1820 ;
      RECT 6.5710 0.7590 8.0210 0.8090 ;
      RECT 7.4990 0.6420 7.5490 0.7590 ;
      RECT 7.1190 0.8090 7.1690 1.2400 ;
      RECT 6.9270 0.5630 6.9770 0.7590 ;
      RECT 6.9270 0.5130 7.1690 0.5630 ;
      RECT 7.1190 0.3830 7.1690 0.5130 ;
      RECT 6.1150 1.5280 10.1510 1.5780 ;
      RECT 6.2670 0.7130 6.5010 0.7630 ;
      RECT 4.7990 0.7670 4.9290 0.8170 ;
      RECT 4.8790 0.5630 4.9290 0.7670 ;
      RECT 4.8390 0.5130 4.9290 0.5630 ;
      RECT 4.7990 0.8170 4.8490 0.9740 ;
      RECT 4.7990 0.9740 4.8890 1.0240 ;
      RECT 4.8390 0.3270 4.8890 0.5130 ;
      RECT 4.8390 1.0240 4.8890 1.1900 ;
      RECT 4.6870 0.2770 4.8890 0.3270 ;
      RECT 4.6870 1.1900 4.8890 1.2400 ;
      RECT 4.6870 0.3270 4.7370 0.5560 ;
      RECT 4.6870 0.9740 4.7370 1.1900 ;
      RECT 5.6590 0.6270 5.9130 0.6770 ;
      RECT 5.8630 0.5630 5.9130 0.6270 ;
      RECT 5.8630 0.6770 5.9130 1.0670 ;
      RECT 5.8630 0.5130 6.7290 0.5630 ;
      RECT 5.8630 1.0670 6.7290 1.1170 ;
      RECT 4.9790 0.4030 5.8010 0.4530 ;
      RECT 5.4470 0.4530 5.4970 0.5770 ;
      RECT 5.7510 0.4530 5.8010 0.5770 ;
      RECT 5.5590 0.4530 5.6090 0.7670 ;
      RECT 5.5590 0.7670 5.8010 0.8170 ;
      RECT 5.7510 0.8170 5.8010 1.2400 ;
      RECT 4.9790 0.4530 5.0290 0.8670 ;
      RECT 4.8990 0.8670 5.0290 0.9170 ;
      RECT 9.8550 0.5620 10.1490 0.6120 ;
      RECT 9.9900 0.4120 10.0400 0.5620 ;
      RECT 9.8550 0.3620 10.0400 0.4120 ;
      RECT 9.8550 0.6120 9.9050 0.8320 ;
      RECT 8.6910 0.8320 9.9050 0.8820 ;
      RECT 9.8550 0.1260 9.9050 0.3620 ;
      RECT 8.6910 0.4200 8.7410 0.8320 ;
      RECT 8.6910 0.3700 8.8590 0.4200 ;
      RECT 1.6870 0.6780 1.9410 0.7020 ;
      RECT 1.6500 0.7020 1.9410 0.7280 ;
      RECT 1.3430 0.4600 1.3930 0.5020 ;
      RECT 1.0230 0.4100 1.3930 0.4600 ;
      RECT 1.3430 0.5020 1.7370 0.5520 ;
      RECT 1.6870 0.5520 1.7370 0.6780 ;
      RECT 1.6500 0.7280 1.7370 0.7520 ;
      RECT 1.6500 0.7520 1.7000 1.0200 ;
      RECT 1.0230 1.0200 1.7000 1.0700 ;
      RECT 2.5590 0.7130 2.6850 0.7630 ;
      RECT 2.5590 0.7630 2.6090 0.8670 ;
      RECT 2.6350 0.5630 2.6850 0.7130 ;
      RECT 2.5590 0.8670 2.8530 0.9170 ;
      RECT 2.5430 0.5130 2.6850 0.5630 ;
      RECT 1.9520 0.9670 3.0050 1.0170 ;
      RECT 1.9520 1.0170 2.0020 1.2140 ;
      RECT 1.9520 0.8280 2.0020 0.9670 ;
      RECT 1.9520 0.7780 2.0410 0.8280 ;
      RECT 1.9910 0.6280 2.0410 0.7780 ;
      RECT 1.9520 0.5780 2.0410 0.6280 ;
      RECT 1.9520 0.3190 2.0020 0.5780 ;
      RECT 5.2950 0.7310 5.3880 0.7810 ;
      RECT 5.2950 0.5050 5.3450 0.7310 ;
      RECT 5.3380 0.7810 5.3880 0.8670 ;
      RECT 5.3380 0.8670 5.5890 0.9170 ;
      RECT 5.3380 0.9170 5.3880 1.0320 ;
      RECT 5.2950 1.0320 5.3880 1.0820 ;
      RECT 5.2950 1.0820 5.3450 1.2400 ;
      RECT 7.9390 1.2000 9.0850 1.2500 ;
      RECT 2.4330 0.4130 2.8370 0.4630 ;
      RECT 2.7870 0.4630 2.8370 0.6800 ;
      RECT 2.4330 0.4630 2.4830 0.6130 ;
      RECT 2.1030 0.6130 2.5490 0.6630 ;
      RECT 2.1030 0.6630 2.1530 0.9120 ;
      RECT 2.1030 0.4130 2.1530 0.6130 ;
      RECT 5.9630 0.6130 6.8650 0.6630 ;
      RECT 6.8150 0.3830 6.8650 0.6130 ;
      RECT 6.1670 0.6630 6.2170 0.9670 ;
      RECT 6.1670 0.9670 6.8650 1.0170 ;
      RECT 6.8150 1.0170 6.8650 1.2400 ;
      RECT 0.7190 0.9410 0.9530 0.9910 ;
      RECT 3.8870 0.8670 4.1690 0.9170 ;
      RECT 4.1190 0.9170 4.1690 1.1270 ;
      RECT 3.0150 1.1270 4.1690 1.1770 ;
      RECT 3.0150 1.1770 3.0650 1.2400 ;
      RECT 3.0150 1.0660 3.1150 1.1270 ;
      RECT 3.0650 0.9170 3.1150 1.0660 ;
      RECT 3.0150 0.4130 3.0650 0.8670 ;
      RECT 3.0150 0.8670 3.3090 0.9170 ;
      RECT 3.8870 0.6070 3.9370 0.8670 ;
      RECT 3.8870 0.5570 3.9770 0.6070 ;
      RECT 3.9270 0.4130 3.9770 0.5570 ;
      RECT 1.1750 1.1330 1.5610 1.1830 ;
      RECT 0.7190 0.5100 1.2570 0.5600 ;
      RECT 0.8870 0.3100 1.5450 0.3600 ;
      RECT 1.4950 0.3600 1.5450 0.3920 ;
      RECT 0.8870 0.3600 0.9370 0.3920 ;
      RECT 3.4710 0.9670 4.0690 1.0170 ;
      RECT 3.1670 0.4070 3.2170 0.6190 ;
      RECT 3.4710 1.0170 3.5210 1.0770 ;
      RECT 3.4710 0.6690 3.5210 0.9670 ;
      RECT 3.1670 0.6190 3.5210 0.6690 ;
      RECT 3.4710 0.4070 3.5210 0.6190 ;
      RECT 4.5950 0.6130 4.8290 0.6630 ;
      RECT 2.4670 1.5240 4.8290 1.5740 ;
      RECT 2.6190 0.0940 4.5250 0.1440 ;
      RECT 4.4430 0.8670 4.6970 0.9170 ;
      RECT 3.3730 1.3900 5.5890 1.4400 ;
      RECT 3.9870 0.6670 4.3730 0.7170 ;
      RECT 7.3990 0.5010 7.7010 0.5510 ;
      RECT 7.6510 0.5510 7.7010 0.6790 ;
      RECT 7.3990 0.5510 7.4490 0.6130 ;
      RECT 7.0270 0.6130 7.4490 0.6630 ;
      RECT 8.4870 1.0620 8.9330 1.1120 ;
      RECT 8.4870 0.1260 8.5370 1.0620 ;
      RECT 1.4520 0.6020 1.6370 0.6520 ;
      RECT 0.2050 0.5260 0.2550 0.8410 ;
      RECT 0.2790 0.8910 0.3290 1.2140 ;
      RECT 0.2050 0.4760 0.3290 0.5260 ;
      RECT 0.2790 0.3160 0.3290 0.4760 ;
      RECT 0.2050 0.8410 1.5020 0.8910 ;
      RECT 1.4520 0.6520 1.5020 0.8410 ;
      RECT 4.5750 0.0920 7.1090 0.1420 ;
      RECT 4.5750 0.1420 4.6250 0.1940 ;
      RECT 4.5350 0.1940 4.6250 0.2440 ;
      RECT 4.5350 0.2440 4.5850 0.5130 ;
      RECT 4.3830 0.5130 4.5850 0.5630 ;
      RECT 4.3830 0.2770 4.4330 0.5130 ;
      RECT 4.4230 0.5630 4.4730 0.7670 ;
      RECT 4.3430 0.7670 4.4730 0.8170 ;
      RECT 4.3430 0.8170 4.3930 0.9670 ;
    LAYER PO ;
      RECT 3.7090 0.0660 3.7390 0.6370 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 2.7970 0.0660 2.8270 0.6910 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 10.7010 0.0660 10.7310 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 4.1650 0.9390 4.1950 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 10.5490 0.0660 10.5790 1.6060 ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 5.9890 0.0660 6.0190 0.6910 ;
      RECT 10.3970 0.0660 10.4270 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 10.0930 0.0660 10.1230 1.6060 ;
      RECT 6.4450 0.0660 6.4750 0.7910 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 10.2450 0.0660 10.2750 1.6060 ;
      RECT 9.7890 0.0660 9.8190 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 4.6210 0.0660 4.6510 0.6910 ;
      RECT 4.1650 0.0660 4.1950 0.6370 ;
      RECT 2.7970 0.8390 2.8270 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 6.4450 0.9390 6.4750 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 4.6210 0.8390 4.6510 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6140 ;
      RECT 9.6370 0.0660 9.6670 1.6060 ;
      RECT 9.3330 0.0660 9.3630 1.6060 ;
      RECT 9.9410 0.0660 9.9710 1.6060 ;
      RECT 5.9890 0.9590 6.0190 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 9.4850 0.0660 9.5150 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 7.9650 0.0670 7.9950 1.6050 ;
      RECT 3.7090 0.9390 3.7390 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
    LAYER NWELL ;
      RECT -0.1150 1.5430 10.9010 1.7870 ;
      RECT -0.1150 0.6790 7.8580 1.5430 ;
      RECT 10.6260 0.6790 10.9010 1.5430 ;
      RECT 8.3200 0.4910 10.1660 1.0830 ;
  END
END RSDFFARX1_LVT

MACRO RSDFFARX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 11.096 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.8790 0.2710 8.5770 0.3210 ;
        RECT 8.4580 0.3210 8.5770 0.3600 ;
        RECT 8.4580 0.2500 8.5770 0.2710 ;
        RECT 7.8790 0.1490 7.9290 0.2710 ;
        RECT 8.5270 0.3600 8.5770 0.9330 ;
        RECT 8.4580 0.2490 8.5690 0.2500 ;
        RECT 7.8790 0.9330 8.5770 0.9830 ;
        RECT 7.8790 0.9830 7.9290 1.2240 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.3040 0.4010 8.4170 0.4020 ;
        RECT 7.5750 0.4020 8.4270 0.4520 ;
        RECT 7.5750 0.1490 7.6250 0.4020 ;
        RECT 8.3040 0.4520 8.4270 0.5120 ;
        RECT 8.3770 0.5120 8.4270 0.8330 ;
        RECT 7.5750 0.8330 8.4270 0.8830 ;
        RECT 7.5750 0.8830 7.6250 1.2240 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 1.1610 1.0110 1.3160 ;
        RECT 0.8890 1.3160 0.9390 1.5240 ;
        RECT 0.8890 1.5240 1.0290 1.5740 ;
    END
    ANTENNAGATEAREA 0.03339 ;
  END D

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6780 0.7250 0.7280 ;
        RECT 0.4010 0.5510 0.5120 0.6780 ;
    END
    ANTENNAGATEAREA 0.06678 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1620 0.0910 1.3330 0.2070 ;
    END
    ANTENNAGATEAREA 0.03339 ;
  END SI

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 8.9270 0.9420 10.3940 1.0020 ;
        RECT 10.2840 0.6900 10.3940 0.9420 ;
    END
  END VDDG

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 11.0960 0.0300 ;
        RECT 2.4070 0.0300 2.4570 0.3070 ;
        RECT 0.4310 0.0300 0.4810 0.4340 ;
        RECT 0.5830 0.0300 0.6330 0.5120 ;
        RECT 1.7990 0.0300 1.8490 0.4050 ;
        RECT 2.2550 0.0300 2.3050 0.5570 ;
        RECT 1.6470 0.0300 1.6970 0.4050 ;
        RECT 8.0310 0.0300 8.0810 0.2210 ;
        RECT 7.7270 0.0300 7.7770 0.3200 ;
        RECT 7.4230 0.0300 7.4730 0.4090 ;
        RECT 10.0070 0.0300 10.0570 0.3120 ;
        RECT 9.7030 0.0300 9.7530 0.2020 ;
        RECT 8.9430 0.0300 8.9930 0.2060 ;
        RECT 7.3110 0.0300 7.3610 0.2830 ;
        RECT 2.4070 0.3070 4.1290 0.3570 ;
        RECT 4.9750 0.2830 7.3610 0.3330 ;
        RECT 3.3190 0.3570 3.3690 0.5580 ;
        RECT 4.0790 0.3570 4.1290 0.5770 ;
        RECT 3.6230 0.3570 3.6730 0.5580 ;
        RECT 7.2710 0.3330 7.3210 0.4430 ;
    END
  END VSS

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0740 1.4650 2.2460 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 11.0960 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 1.7990 1.1310 1.8490 1.6420 ;
        RECT 1.6470 1.1310 1.6970 1.6420 ;
        RECT 2.3670 1.3400 2.4170 1.6420 ;
        RECT 5.6390 1.3400 5.6890 1.6420 ;
        RECT 2.2370 1.2900 8.0810 1.3400 ;
        RECT 4.9910 0.9730 5.0410 1.2900 ;
        RECT 8.0310 1.0530 8.0810 1.2900 ;
        RECT 7.7270 0.9610 7.7770 1.2900 ;
        RECT 7.4230 0.9130 7.4730 1.2900 ;
    END
  END VDD

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.1140 0.8510 5.2680 0.9670 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END RSTB

  PIN RETN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.9450 1.4080 9.6340 1.4580 ;
        RECT 9.5220 1.3130 9.6340 1.4080 ;
    END
    ANTENNAGATEAREA 0.084 ;
  END RETN
  OBS
    LAYER M1 ;
      RECT 4.3830 0.2770 4.4330 0.5130 ;
      RECT 4.4230 0.5630 4.4730 0.7670 ;
      RECT 4.3430 0.7670 4.4730 0.8170 ;
      RECT 4.3430 0.8170 4.3930 0.9670 ;
      RECT 4.3430 0.9670 4.4330 1.0170 ;
      RECT 4.3830 1.0170 4.4330 1.1900 ;
      RECT 4.3830 1.1900 4.5850 1.2400 ;
      RECT 4.5350 0.9740 4.5850 1.1900 ;
      RECT 6.1150 1.5280 10.4550 1.5780 ;
      RECT 1.4520 0.6020 1.6370 0.6520 ;
      RECT 0.2050 0.8410 1.5020 0.8910 ;
      RECT 1.4520 0.6520 1.5020 0.8410 ;
      RECT 0.2050 0.5260 0.2550 0.8410 ;
      RECT 0.2790 0.8910 0.3290 1.2140 ;
      RECT 0.2050 0.4760 0.3290 0.5260 ;
      RECT 0.2790 0.3160 0.3290 0.4760 ;
      RECT 1.6870 0.6780 1.9410 0.7020 ;
      RECT 1.6500 0.7020 1.9410 0.7280 ;
      RECT 1.0230 0.4100 1.3930 0.4600 ;
      RECT 1.3430 0.4600 1.3930 0.5020 ;
      RECT 1.3430 0.5020 1.7370 0.5520 ;
      RECT 1.6870 0.5520 1.7370 0.6780 ;
      RECT 1.6500 0.7280 1.7370 0.7520 ;
      RECT 1.6500 0.7520 1.7000 1.0200 ;
      RECT 1.0230 1.0200 1.7000 1.0700 ;
      RECT 0.7190 0.5100 1.2570 0.5600 ;
      RECT 0.8870 0.3100 1.5450 0.3600 ;
      RECT 0.8870 0.3600 0.9370 0.3920 ;
      RECT 1.4950 0.3600 1.5450 0.3920 ;
      RECT 1.9520 0.9670 3.0050 1.0170 ;
      RECT 1.9520 1.0170 2.0020 1.2140 ;
      RECT 1.9520 0.8280 2.0020 0.9670 ;
      RECT 1.9520 0.7780 2.0410 0.8280 ;
      RECT 1.9910 0.6280 2.0410 0.7780 ;
      RECT 1.9520 0.5780 2.0410 0.6280 ;
      RECT 1.9520 0.3190 2.0020 0.5780 ;
      RECT 2.5430 0.5130 2.6850 0.5630 ;
      RECT 2.6350 0.5630 2.6850 0.7130 ;
      RECT 2.5590 0.7130 2.6850 0.7630 ;
      RECT 2.5590 0.7630 2.6090 0.8670 ;
      RECT 2.5590 0.8670 2.8530 0.9170 ;
      RECT 2.1030 0.6130 2.5490 0.6630 ;
      RECT 2.4330 0.4630 2.4830 0.6130 ;
      RECT 2.4330 0.4130 2.8370 0.4630 ;
      RECT 2.7870 0.4630 2.8370 0.6800 ;
      RECT 2.1030 0.6630 2.1530 0.9120 ;
      RECT 2.1030 0.4130 2.1530 0.6130 ;
      RECT 3.8870 0.8670 4.1690 0.9170 ;
      RECT 4.1190 0.9170 4.1690 1.1270 ;
      RECT 3.0150 1.1270 4.1690 1.1770 ;
      RECT 3.0150 1.1770 3.0650 1.2400 ;
      RECT 3.0150 1.0660 3.1150 1.1270 ;
      RECT 3.0650 0.9170 3.1150 1.0660 ;
      RECT 3.0150 0.4130 3.0650 0.8670 ;
      RECT 3.0150 0.8670 3.3090 0.9170 ;
      RECT 3.8870 0.6070 3.9370 0.8670 ;
      RECT 3.8870 0.5570 3.9770 0.6070 ;
      RECT 3.9270 0.4130 3.9770 0.5570 ;
      RECT 3.4710 0.9670 4.0690 1.0170 ;
      RECT 3.1670 0.4070 3.2170 0.6190 ;
      RECT 3.4710 1.0170 3.5210 1.0770 ;
      RECT 3.4710 0.6690 3.5210 0.9670 ;
      RECT 3.1670 0.6190 3.5210 0.6690 ;
      RECT 3.4710 0.4070 3.5210 0.6190 ;
      RECT 2.6190 0.0940 4.5250 0.1440 ;
      RECT 5.8630 0.5130 6.7290 0.5630 ;
      RECT 5.8630 0.5630 5.9130 0.6270 ;
      RECT 5.6590 0.6270 5.9130 0.6770 ;
      RECT 5.8630 0.6770 5.9130 1.0670 ;
      RECT 5.8630 1.0670 6.7290 1.1170 ;
      RECT 4.9790 0.4030 5.8010 0.4530 ;
      RECT 5.4470 0.4530 5.4970 0.5770 ;
      RECT 5.7510 0.4530 5.8010 0.5770 ;
      RECT 5.5590 0.4530 5.6090 0.7670 ;
      RECT 5.5590 0.7670 5.8010 0.8170 ;
      RECT 5.7510 0.8170 5.8010 1.2400 ;
      RECT 4.9790 0.4530 5.0290 0.8670 ;
      RECT 4.8990 0.8670 5.0290 0.9170 ;
      RECT 4.8390 0.5130 4.9290 0.5630 ;
      RECT 4.8790 0.5630 4.9290 0.7670 ;
      RECT 4.7990 0.7670 4.9290 0.8170 ;
      RECT 4.6870 0.2770 4.8890 0.3270 ;
      RECT 4.6870 0.3270 4.7370 0.5560 ;
      RECT 4.8390 0.3270 4.8890 0.5130 ;
      RECT 4.7990 0.8170 4.8490 0.9740 ;
      RECT 4.7990 0.9740 4.8890 1.0240 ;
      RECT 4.8390 1.0240 4.8890 1.1900 ;
      RECT 4.6870 1.1900 4.8890 1.2400 ;
      RECT 4.6870 0.9740 4.7370 1.1900 ;
      RECT 5.2950 0.7310 5.3880 0.7810 ;
      RECT 5.2950 0.5050 5.3450 0.7310 ;
      RECT 5.3380 0.7810 5.3880 0.8670 ;
      RECT 5.3380 0.8670 5.5890 0.9170 ;
      RECT 5.3380 0.9170 5.3880 1.0320 ;
      RECT 5.2950 1.0320 5.3880 1.0820 ;
      RECT 5.2950 1.0820 5.3450 1.2400 ;
      RECT 6.5710 0.7130 8.3250 0.7630 ;
      RECT 7.1190 0.7630 7.1690 1.2400 ;
      RECT 6.9270 0.5630 6.9770 0.7130 ;
      RECT 6.9270 0.5130 7.1690 0.5630 ;
      RECT 7.1190 0.3830 7.1690 0.5130 ;
      RECT 7.4990 0.6420 7.5490 0.7130 ;
      RECT 7.6510 0.6420 7.7010 0.7130 ;
      RECT 7.0270 0.6130 7.4010 0.6630 ;
      RECT 7.3500 0.5700 7.4010 0.6130 ;
      RECT 7.3500 0.5200 7.8350 0.5700 ;
      RECT 7.7850 0.5700 7.8350 0.6040 ;
      RECT 7.7850 0.6040 8.0210 0.6540 ;
      RECT 5.9630 0.6130 6.8650 0.6630 ;
      RECT 6.8150 0.3830 6.8650 0.6130 ;
      RECT 6.1670 0.6630 6.2170 0.9670 ;
      RECT 6.1670 0.9670 6.8650 1.0170 ;
      RECT 6.8150 1.0170 6.8650 1.2400 ;
      RECT 8.7910 1.0620 9.2370 1.1120 ;
      RECT 8.7910 0.1260 8.8410 1.0620 ;
      RECT 9.5510 0.4620 9.8450 0.5120 ;
      RECT 9.5510 0.1820 9.6010 0.4620 ;
      RECT 9.5510 0.5120 9.6010 0.6350 ;
      RECT 9.2310 0.1320 9.6010 0.1820 ;
      RECT 9.2310 0.6350 9.6010 0.6850 ;
      RECT 9.8550 0.5890 10.0480 0.6390 ;
      RECT 9.9980 0.5120 10.0480 0.5890 ;
      RECT 9.9980 0.4620 10.1490 0.5120 ;
      RECT 9.9980 0.4120 10.0480 0.4620 ;
      RECT 9.8550 0.3620 10.0480 0.4120 ;
      RECT 9.8550 0.6390 9.9050 0.7820 ;
      RECT 9.8550 0.1260 9.9050 0.3620 ;
      RECT 9.0950 0.4940 9.4490 0.5440 ;
      RECT 9.3990 0.3480 9.4490 0.4940 ;
      RECT 9.0950 0.5440 9.1450 0.7820 ;
      RECT 10.1590 0.5620 10.4530 0.6120 ;
      RECT 10.2940 0.4120 10.3440 0.5620 ;
      RECT 10.1590 0.3620 10.3440 0.4120 ;
      RECT 10.1590 0.6120 10.2090 0.8320 ;
      RECT 8.9950 0.8320 10.2090 0.8820 ;
      RECT 10.1590 0.1260 10.2090 0.3620 ;
      RECT 8.9950 0.4200 9.0450 0.8320 ;
      RECT 8.9950 0.3700 9.1630 0.4200 ;
      RECT 0.7190 0.9410 0.9530 0.9910 ;
      RECT 3.3730 1.3900 5.5890 1.4400 ;
      RECT 1.1750 1.1330 1.5610 1.1830 ;
      RECT 2.4670 1.5240 4.8290 1.5740 ;
      RECT 3.9870 0.6670 4.3730 0.7170 ;
      RECT 4.5950 0.6130 4.8290 0.6630 ;
      RECT 4.4430 0.8670 4.6970 0.9170 ;
      RECT 6.2670 0.7130 6.5010 0.7630 ;
      RECT 8.2430 1.2000 9.3890 1.2500 ;
      RECT 4.5750 0.0920 7.1090 0.1420 ;
      RECT 4.5750 0.1420 4.6250 0.1940 ;
      RECT 4.5350 0.1940 4.6250 0.2440 ;
      RECT 4.5350 0.2440 4.5850 0.5130 ;
      RECT 4.3830 0.5130 4.5850 0.5630 ;
    LAYER PO ;
      RECT 9.9410 0.0660 9.9710 1.6060 ;
      RECT 9.6370 0.0660 9.6670 1.6060 ;
      RECT 10.2450 0.0660 10.2750 1.6060 ;
      RECT 5.9890 0.9590 6.0190 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 9.7890 0.0660 9.8190 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 8.2690 0.0670 8.2990 1.6050 ;
      RECT 3.7090 0.9390 3.7390 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
      RECT 3.7090 0.0660 3.7390 0.6370 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 2.7970 0.0660 2.8270 0.6910 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 11.0050 0.0660 11.0350 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 4.1650 0.9390 4.1950 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 10.8530 0.0660 10.8830 1.6060 ;
      RECT 9.4850 0.0660 9.5150 1.6060 ;
      RECT 5.9890 0.0660 6.0190 0.6910 ;
      RECT 10.7010 0.0660 10.7310 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 10.3970 0.0660 10.4270 1.6060 ;
      RECT 6.4450 0.0660 6.4750 0.7910 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 10.5490 0.0660 10.5790 1.6060 ;
      RECT 10.0930 0.0660 10.1230 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 4.6210 0.0660 4.6510 0.6910 ;
      RECT 4.1650 0.0660 4.1950 0.6370 ;
      RECT 2.7970 0.8390 2.8270 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 6.4450 0.9390 6.4750 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 4.6210 0.8390 4.6510 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 9.3330 0.0660 9.3630 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6140 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
    LAYER NWELL ;
      RECT -0.1160 1.5430 11.2040 1.7730 ;
      RECT -0.1160 0.6790 8.1620 1.5430 ;
      RECT 10.9290 0.6790 11.2040 1.5430 ;
      RECT 8.6230 0.4910 10.4690 1.0830 ;
  END
END RSDFFARX2_LVT

MACRO RSDFFNARX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.792 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 1.1610 1.0110 1.3160 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6780 0.7250 0.7280 ;
        RECT 0.4010 0.5510 0.5120 0.6780 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1620 0.0970 1.3180 0.2070 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 8.6230 0.9420 10.0900 1.0020 ;
        RECT 9.9800 0.6900 10.0900 0.9420 ;
    END
  END VDDG

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 10.7920 0.0300 ;
        RECT 9.7030 0.0300 9.7530 0.3120 ;
        RECT 1.7990 0.0300 1.8490 0.4050 ;
        RECT 9.3990 0.0300 9.4490 0.2020 ;
        RECT 0.4310 0.0300 0.4810 0.4340 ;
        RECT 0.5830 0.0300 0.6330 0.5120 ;
        RECT 8.6390 0.0300 8.6890 0.2060 ;
        RECT 7.5750 0.0300 7.6250 0.2410 ;
        RECT 1.6470 0.0300 1.6970 0.4050 ;
        RECT 2.2090 0.0300 2.2590 0.3070 ;
        RECT 7.3110 0.0300 7.3610 0.2830 ;
        RECT 2.2090 0.3070 4.1290 0.3570 ;
        RECT 4.9750 0.2830 7.3610 0.3330 ;
        RECT 2.2550 0.3570 2.3050 0.5570 ;
        RECT 4.0790 0.3570 4.1290 0.5770 ;
        RECT 3.3190 0.3570 3.3690 0.5580 ;
        RECT 3.6230 0.3570 3.6730 0.5580 ;
        RECT 7.2710 0.3330 7.3210 0.4430 ;
    END
  END VSS

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0740 1.4650 2.2460 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.7270 0.9690 8.2610 1.0190 ;
        RECT 7.7270 1.0190 7.9610 1.1290 ;
        RECT 8.2110 0.3510 8.2610 0.9690 ;
        RECT 7.7270 1.1290 7.7770 1.3270 ;
        RECT 7.7110 0.3010 8.2610 0.3510 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.4230 0.1570 7.4730 0.4010 ;
        RECT 7.4230 0.4010 8.1230 0.4510 ;
        RECT 8.0010 0.4510 8.1230 0.5380 ;
        RECT 8.0730 0.5380 8.1230 0.8590 ;
        RECT 7.4230 0.8590 8.1230 0.9090 ;
        RECT 7.4230 0.9090 7.4730 1.2320 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 10.7920 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 1.7990 1.1310 1.8490 1.6420 ;
        RECT 1.6470 1.1310 1.6970 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 5.6390 1.3400 5.6890 1.6420 ;
        RECT 2.3670 1.3400 2.4170 1.6420 ;
        RECT 2.2370 1.2900 7.6250 1.3400 ;
        RECT 7.5750 0.9590 7.6250 1.2900 ;
        RECT 4.9910 0.9730 5.0410 1.2900 ;
    END
  END VDD

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.1140 0.8510 5.2680 0.9670 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END RSTB

  PIN RETN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.9450 1.4080 9.3300 1.4580 ;
        RECT 9.2180 1.3130 9.3300 1.4080 ;
    END
    ANTENNAGATEAREA 0.084 ;
  END RETN
  OBS
    LAYER M1 ;
      RECT 4.3830 1.1900 4.5850 1.2400 ;
      RECT 4.5350 0.9740 4.5850 1.1900 ;
      RECT 8.7910 0.4940 9.1450 0.5440 ;
      RECT 8.7910 0.5440 8.8410 0.7820 ;
      RECT 9.0950 0.3480 9.1450 0.4940 ;
      RECT 9.2470 0.4620 9.5410 0.5120 ;
      RECT 9.2470 0.5120 9.2970 0.6350 ;
      RECT 9.2470 0.1820 9.2970 0.4620 ;
      RECT 8.9270 0.6350 9.2970 0.6850 ;
      RECT 8.9270 0.1320 9.2970 0.1820 ;
      RECT 6.5710 0.7590 8.0210 0.8090 ;
      RECT 7.4990 0.6420 7.5490 0.7590 ;
      RECT 7.1190 0.8090 7.1690 1.2400 ;
      RECT 6.9270 0.5630 6.9770 0.7590 ;
      RECT 6.9270 0.5130 7.1690 0.5630 ;
      RECT 7.1190 0.3830 7.1690 0.5130 ;
      RECT 6.1150 1.5280 10.1510 1.5780 ;
      RECT 6.2670 0.7130 6.5010 0.7630 ;
      RECT 9.6940 0.4120 9.7440 0.4620 ;
      RECT 9.6940 0.4620 9.8450 0.5120 ;
      RECT 9.6940 0.5120 9.7440 0.5890 ;
      RECT 9.5510 0.5890 9.7440 0.6390 ;
      RECT 9.5510 0.3620 9.7440 0.4120 ;
      RECT 9.5510 0.1260 9.6010 0.3620 ;
      RECT 9.5510 0.6390 9.6010 0.7820 ;
      RECT 4.7990 0.7670 4.9290 0.8170 ;
      RECT 4.8790 0.5630 4.9290 0.7670 ;
      RECT 4.8390 0.5130 4.9290 0.5630 ;
      RECT 4.6870 1.1900 4.8890 1.2400 ;
      RECT 4.6870 0.9740 4.7370 1.1900 ;
      RECT 4.8390 1.0240 4.8890 1.1900 ;
      RECT 4.7990 0.9740 4.8890 1.0240 ;
      RECT 4.7990 0.8170 4.8490 0.9740 ;
      RECT 4.8390 0.3270 4.8890 0.5130 ;
      RECT 4.6870 0.2770 4.8890 0.3270 ;
      RECT 4.6870 0.3270 4.7370 0.5560 ;
      RECT 5.6590 0.6270 5.9130 0.6770 ;
      RECT 5.8630 0.5630 5.9130 0.6270 ;
      RECT 5.8630 0.6770 5.9130 1.0670 ;
      RECT 5.8630 0.5130 6.7290 0.5630 ;
      RECT 5.8630 1.0670 6.7290 1.1170 ;
      RECT 4.9790 0.4030 5.8010 0.4530 ;
      RECT 5.4470 0.4530 5.4970 0.5770 ;
      RECT 5.7510 0.4530 5.8010 0.5770 ;
      RECT 5.5590 0.4530 5.6090 0.7670 ;
      RECT 5.5590 0.7670 5.8010 0.8170 ;
      RECT 5.7510 0.8170 5.8010 1.2400 ;
      RECT 4.9790 0.4530 5.0290 0.8670 ;
      RECT 4.8990 0.8670 5.0290 0.9170 ;
      RECT 9.8550 0.5620 10.1490 0.6120 ;
      RECT 9.9900 0.4120 10.0400 0.5620 ;
      RECT 9.8550 0.3620 10.0400 0.4120 ;
      RECT 9.8550 0.6120 9.9050 0.8320 ;
      RECT 8.6910 0.8320 9.9050 0.8820 ;
      RECT 9.8550 0.1260 9.9050 0.3620 ;
      RECT 8.6910 0.4200 8.7410 0.8320 ;
      RECT 8.6910 0.3700 8.8590 0.4200 ;
      RECT 1.6870 0.6780 1.9410 0.7020 ;
      RECT 1.6500 0.7020 1.9410 0.7280 ;
      RECT 1.3430 0.4600 1.3930 0.5020 ;
      RECT 1.0230 0.4100 1.3930 0.4600 ;
      RECT 1.3430 0.5020 1.7370 0.5520 ;
      RECT 1.6870 0.5520 1.7370 0.6780 ;
      RECT 1.6500 0.7280 1.7370 0.7520 ;
      RECT 1.6500 0.7520 1.7000 1.0200 ;
      RECT 1.0230 1.0200 1.7000 1.0700 ;
      RECT 1.9520 0.9670 3.0050 1.0170 ;
      RECT 1.9520 1.0170 2.0020 1.2140 ;
      RECT 1.9520 0.8280 2.0020 0.9670 ;
      RECT 1.9520 0.7780 2.0410 0.8280 ;
      RECT 1.9910 0.6280 2.0410 0.7780 ;
      RECT 1.9520 0.5780 2.0410 0.6280 ;
      RECT 1.9520 0.3190 2.0020 0.5780 ;
      RECT 5.2950 0.7310 5.3880 0.7810 ;
      RECT 5.2950 0.5050 5.3450 0.7310 ;
      RECT 5.3380 0.7810 5.3880 0.8670 ;
      RECT 5.3380 0.8670 5.5890 0.9170 ;
      RECT 5.3380 0.9170 5.3880 1.0320 ;
      RECT 5.2950 1.0320 5.3880 1.0820 ;
      RECT 5.2950 1.0820 5.3450 1.2400 ;
      RECT 7.9390 1.2000 9.0850 1.2500 ;
      RECT 5.9630 0.6130 6.8650 0.6630 ;
      RECT 6.8150 0.3830 6.8650 0.6130 ;
      RECT 6.1670 0.6630 6.2170 0.9670 ;
      RECT 6.1670 0.9670 6.8650 1.0170 ;
      RECT 6.8150 1.0170 6.8650 1.2400 ;
      RECT 0.7190 0.9410 0.9530 0.9910 ;
      RECT 3.8870 0.8670 4.1690 0.9170 ;
      RECT 4.1190 0.9170 4.1690 1.1270 ;
      RECT 3.0150 1.1270 4.1690 1.1770 ;
      RECT 3.0150 1.1770 3.0650 1.2400 ;
      RECT 3.0150 1.0660 3.1150 1.1270 ;
      RECT 3.0650 0.9170 3.1150 1.0660 ;
      RECT 3.0150 0.4130 3.0650 0.8670 ;
      RECT 3.0150 0.8670 3.3090 0.9170 ;
      RECT 3.8870 0.6070 3.9370 0.8670 ;
      RECT 3.8870 0.5570 3.9770 0.6070 ;
      RECT 3.9270 0.4130 3.9770 0.5570 ;
      RECT 2.5430 0.5130 2.6850 0.5630 ;
      RECT 2.6350 0.5630 2.6850 0.6130 ;
      RECT 2.6350 0.6130 2.8680 0.6630 ;
      RECT 2.6350 0.6630 2.6850 0.7540 ;
      RECT 2.5420 0.7540 2.6850 0.8040 ;
      RECT 1.1750 1.1330 1.5610 1.1830 ;
      RECT 0.7190 0.5100 1.2570 0.5600 ;
      RECT 0.8870 0.3100 1.5450 0.3600 ;
      RECT 1.4950 0.3600 1.5450 0.3920 ;
      RECT 0.8870 0.3600 0.9370 0.3920 ;
      RECT 3.4710 0.9670 4.0690 1.0170 ;
      RECT 3.1670 0.4070 3.2170 0.6190 ;
      RECT 3.4710 1.0170 3.5210 1.0770 ;
      RECT 3.4710 0.6690 3.5210 0.9670 ;
      RECT 3.1670 0.6190 3.5210 0.6690 ;
      RECT 3.4710 0.4070 3.5210 0.6190 ;
      RECT 4.5950 0.6130 4.8290 0.6630 ;
      RECT 2.6190 1.5240 4.8290 1.5740 ;
      RECT 2.3150 0.0940 4.5250 0.1440 ;
      RECT 4.4430 0.8670 4.6970 0.9170 ;
      RECT 2.1030 0.6130 2.5490 0.6630 ;
      RECT 2.1030 0.8670 2.8530 0.9170 ;
      RECT 2.1030 0.4130 2.1530 0.6130 ;
      RECT 2.1030 0.6630 2.1530 0.8670 ;
      RECT 3.3730 1.3900 5.5890 1.4400 ;
      RECT 3.9870 0.6670 4.3730 0.7170 ;
      RECT 7.3990 0.5010 7.7010 0.5510 ;
      RECT 7.6510 0.5510 7.7010 0.6790 ;
      RECT 7.3990 0.5510 7.4490 0.6130 ;
      RECT 7.0270 0.6130 7.4490 0.6630 ;
      RECT 8.4870 1.0620 8.9330 1.1120 ;
      RECT 8.4870 0.1260 8.5370 1.0620 ;
      RECT 1.4520 0.6020 1.6370 0.6520 ;
      RECT 0.2050 0.5260 0.2550 0.8410 ;
      RECT 0.2790 0.8910 0.3290 1.2140 ;
      RECT 0.2050 0.4760 0.3290 0.5260 ;
      RECT 0.2790 0.3160 0.3290 0.4760 ;
      RECT 0.2050 0.8410 1.5020 0.8910 ;
      RECT 1.4520 0.6520 1.5020 0.8410 ;
      RECT 4.5750 0.0920 7.1090 0.1420 ;
      RECT 4.5750 0.1420 4.6250 0.1940 ;
      RECT 4.5350 0.1940 4.6250 0.2440 ;
      RECT 4.5350 0.2440 4.5850 0.5130 ;
      RECT 4.3830 0.5130 4.5850 0.5630 ;
      RECT 4.3830 0.2770 4.4330 0.5130 ;
      RECT 4.4230 0.5630 4.4730 0.7670 ;
      RECT 4.3430 0.7670 4.4730 0.8170 ;
      RECT 4.3430 0.8170 4.3930 0.9670 ;
      RECT 4.3430 0.9670 4.4330 1.0170 ;
      RECT 4.3830 1.0170 4.4330 1.1900 ;
    LAYER PO ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 2.7970 0.0660 2.8270 0.6910 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 10.7010 0.0660 10.7310 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 4.1650 0.9390 4.1950 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 10.5490 0.0660 10.5790 1.6060 ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 5.9890 0.0660 6.0190 0.6910 ;
      RECT 10.3970 0.0660 10.4270 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 10.0930 0.0660 10.1230 1.6060 ;
      RECT 6.4450 0.0660 6.4750 0.7910 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 10.2450 0.0660 10.2750 1.6060 ;
      RECT 9.7890 0.0660 9.8190 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 4.6210 0.0660 4.6510 0.6910 ;
      RECT 4.1650 0.0660 4.1950 0.6370 ;
      RECT 2.7970 0.8390 2.8270 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 6.4450 0.9390 6.4750 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 4.6210 0.8390 4.6510 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6140 ;
      RECT 9.6370 0.0660 9.6670 1.6060 ;
      RECT 9.3330 0.0660 9.3630 1.6060 ;
      RECT 9.9410 0.0660 9.9710 1.6060 ;
      RECT 5.9890 0.9590 6.0190 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 9.4850 0.0660 9.5150 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 7.9650 0.0670 7.9950 1.6050 ;
      RECT 3.7090 0.9390 3.7390 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
      RECT 3.7090 0.0660 3.7390 0.6370 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
    LAYER NWELL ;
      RECT -0.1160 1.5430 10.9000 1.7730 ;
      RECT -0.1160 0.6790 7.8580 1.5430 ;
      RECT 10.6250 0.6790 10.9000 1.5430 ;
      RECT 8.3190 0.4910 10.1650 1.0830 ;
  END
END RSDFFNARX1_LVT

MACRO RSDFFNARX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 11.096 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 1.1610 1.0110 1.3160 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6780 0.7250 0.7280 ;
        RECT 0.4010 0.5510 0.5120 0.6780 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1620 0.0970 1.3180 0.2070 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.8790 0.2710 8.5770 0.3210 ;
        RECT 8.4590 0.3210 8.5770 0.3590 ;
        RECT 8.4590 0.2500 8.5770 0.2710 ;
        RECT 7.8790 0.1490 7.9290 0.2710 ;
        RECT 8.5270 0.3590 8.5770 0.9330 ;
        RECT 8.4590 0.2490 8.5690 0.2500 ;
        RECT 7.8790 0.9330 8.5770 0.9830 ;
        RECT 7.8790 0.9830 7.9290 1.2240 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 8.9270 0.9420 10.3940 1.0020 ;
        RECT 10.2840 0.6900 10.3940 0.9420 ;
    END
  END VDDG

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.3050 0.4010 8.4170 0.4020 ;
        RECT 7.5750 0.4020 8.4270 0.4520 ;
        RECT 7.5750 0.1490 7.6250 0.4020 ;
        RECT 8.3050 0.4520 8.4270 0.5120 ;
        RECT 8.3770 0.5120 8.4270 0.8330 ;
        RECT 7.5750 0.8330 8.4270 0.8830 ;
        RECT 7.5750 0.8830 7.6250 1.2240 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 11.0960 0.0300 ;
        RECT 10.0060 0.0300 10.0560 0.3120 ;
        RECT 1.7980 0.0300 1.8480 0.4050 ;
        RECT 8.0300 0.0300 8.0800 0.2210 ;
        RECT 9.7020 0.0300 9.7520 0.2020 ;
        RECT 0.4300 0.0300 0.4800 0.4340 ;
        RECT 0.5820 0.0300 0.6320 0.5120 ;
        RECT 8.9420 0.0300 8.9920 0.2060 ;
        RECT 7.4220 0.0300 7.4720 0.4090 ;
        RECT 1.6460 0.0300 1.6960 0.4050 ;
        RECT 7.7260 0.0300 7.7760 0.3200 ;
        RECT 7.3100 0.0300 7.3600 0.2830 ;
        RECT 2.2090 0.0300 2.2590 0.3070 ;
        RECT 4.9750 0.2830 7.3610 0.3330 ;
        RECT 2.2090 0.3070 4.1290 0.3570 ;
        RECT 7.2710 0.3330 7.3210 0.4430 ;
        RECT 2.2550 0.3570 2.3050 0.5570 ;
        RECT 4.0790 0.3570 4.1290 0.5770 ;
        RECT 3.3190 0.3570 3.3690 0.5580 ;
        RECT 3.6230 0.3570 3.6730 0.5580 ;
    END
  END VSS

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0740 1.4650 2.2460 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 11.0960 1.7020 ;
        RECT 0.5820 1.0330 0.6320 1.6420 ;
        RECT 1.7980 1.1310 1.8480 1.6420 ;
        RECT 1.6460 1.1310 1.6960 1.6420 ;
        RECT 0.4300 1.0330 0.4800 1.6420 ;
        RECT 2.3660 1.3400 2.4160 1.6420 ;
        RECT 5.6530 1.3400 5.7030 1.6420 ;
        RECT 2.2370 1.2900 8.0810 1.3400 ;
        RECT 8.0310 1.0530 8.0810 1.2900 ;
        RECT 7.4230 0.9130 7.4730 1.2900 ;
        RECT 7.7270 0.9610 7.7770 1.2900 ;
        RECT 4.9910 0.9730 5.0410 1.2900 ;
    END
  END VDD

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.1140 0.8510 5.2680 0.9670 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END RSTB

  PIN RETN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.9450 1.4080 9.6340 1.4580 ;
        RECT 9.5220 1.3130 9.6340 1.4080 ;
    END
    ANTENNAGATEAREA 0.084 ;
  END RETN
  OBS
    LAYER M1 ;
      RECT 1.4520 0.6520 1.5020 0.8410 ;
      RECT 4.5750 0.0920 7.1090 0.1420 ;
      RECT 4.5750 0.1420 4.6250 0.1940 ;
      RECT 4.5350 0.1940 4.6250 0.2440 ;
      RECT 4.5350 0.2440 4.5850 0.5130 ;
      RECT 4.3830 0.5130 4.5850 0.5630 ;
      RECT 4.3830 0.2770 4.4330 0.5130 ;
      RECT 4.4230 0.5630 4.4730 0.7670 ;
      RECT 4.3430 0.7670 4.4730 0.8170 ;
      RECT 4.3430 0.8170 4.3930 0.9670 ;
      RECT 4.3430 0.9670 4.4330 1.0170 ;
      RECT 4.3830 1.0170 4.4330 1.1900 ;
      RECT 4.3830 1.1900 4.5850 1.2400 ;
      RECT 4.5350 0.9740 4.5850 1.1900 ;
      RECT 5.9630 0.6130 6.8650 0.6630 ;
      RECT 6.8150 0.3830 6.8650 0.6130 ;
      RECT 6.1670 0.6630 6.2170 0.9670 ;
      RECT 6.1670 0.9670 6.8650 1.0170 ;
      RECT 6.8150 1.0170 6.8650 1.2400 ;
      RECT 4.9790 0.4030 5.8010 0.4530 ;
      RECT 5.4470 0.4530 5.4970 0.5770 ;
      RECT 5.7510 0.4530 5.8010 0.5770 ;
      RECT 5.5590 0.4530 5.6090 0.7670 ;
      RECT 5.5590 0.7670 5.8010 0.8170 ;
      RECT 5.7510 0.8170 5.8010 1.2400 ;
      RECT 4.9790 0.4530 5.0290 0.8670 ;
      RECT 4.8990 0.8670 5.0290 0.9170 ;
      RECT 9.5510 0.4620 9.8450 0.5120 ;
      RECT 9.5510 0.1820 9.6010 0.4620 ;
      RECT 9.2310 0.1320 9.6010 0.1820 ;
      RECT 9.5510 0.5120 9.6010 0.6350 ;
      RECT 9.2310 0.6350 9.6010 0.6850 ;
      RECT 9.8550 0.5890 10.0480 0.6390 ;
      RECT 9.9980 0.5120 10.0480 0.5890 ;
      RECT 9.9980 0.4620 10.1490 0.5120 ;
      RECT 9.9980 0.4120 10.0480 0.4620 ;
      RECT 9.8550 0.3620 10.0480 0.4120 ;
      RECT 9.8550 0.6390 9.9050 0.7820 ;
      RECT 9.8550 0.1260 9.9050 0.3620 ;
      RECT 1.9520 0.9670 3.0050 1.0170 ;
      RECT 1.9520 1.0170 2.0020 1.2140 ;
      RECT 1.9520 0.8280 2.0020 0.9670 ;
      RECT 1.9520 0.7780 2.0410 0.8280 ;
      RECT 1.9910 0.6280 2.0410 0.7780 ;
      RECT 1.9520 0.5780 2.0410 0.6280 ;
      RECT 1.9520 0.3190 2.0020 0.5780 ;
      RECT 9.0950 0.4940 9.4490 0.5440 ;
      RECT 9.3990 0.3480 9.4490 0.4940 ;
      RECT 9.0950 0.5440 9.1450 0.7820 ;
      RECT 6.5710 0.7210 8.3250 0.7710 ;
      RECT 7.1190 0.7710 7.1690 1.2400 ;
      RECT 6.9270 0.5630 6.9770 0.7210 ;
      RECT 6.9270 0.5130 7.1690 0.5630 ;
      RECT 7.1190 0.3830 7.1690 0.5130 ;
      RECT 7.4990 0.6420 7.5490 0.7210 ;
      RECT 7.6510 0.6420 7.7010 0.7210 ;
      RECT 6.1150 1.5280 10.4550 1.5780 ;
      RECT 6.2670 0.7130 6.5010 0.7630 ;
      RECT 4.8390 0.5130 4.9290 0.5630 ;
      RECT 4.8790 0.5630 4.9290 0.7670 ;
      RECT 4.7990 0.7670 4.9290 0.8170 ;
      RECT 4.6870 0.2770 4.8890 0.3270 ;
      RECT 4.6870 0.3270 4.7370 0.5560 ;
      RECT 4.8390 0.3270 4.8890 0.5130 ;
      RECT 4.7990 0.8170 4.8490 0.9740 ;
      RECT 4.7990 0.9740 4.8890 1.0240 ;
      RECT 4.8390 1.0240 4.8890 1.1900 ;
      RECT 4.6870 1.1900 4.8890 1.2400 ;
      RECT 4.6870 0.9740 4.7370 1.1900 ;
      RECT 5.6590 0.6270 5.9130 0.6770 ;
      RECT 5.8630 0.5630 5.9130 0.6270 ;
      RECT 5.8630 0.6770 5.9130 1.0670 ;
      RECT 5.8630 0.5130 6.7290 0.5630 ;
      RECT 5.8630 1.0670 6.7290 1.1170 ;
      RECT 10.1590 0.5620 10.4530 0.6120 ;
      RECT 10.2940 0.4120 10.3440 0.5620 ;
      RECT 10.1590 0.3620 10.3440 0.4120 ;
      RECT 10.1590 0.6120 10.2090 0.8320 ;
      RECT 8.9950 0.8320 10.2090 0.8820 ;
      RECT 10.1590 0.1260 10.2090 0.3620 ;
      RECT 8.9950 0.4200 9.0450 0.8320 ;
      RECT 8.9950 0.3700 9.1630 0.4200 ;
      RECT 1.6870 0.6780 1.9410 0.7020 ;
      RECT 1.6500 0.7020 1.9410 0.7280 ;
      RECT 1.3430 0.4600 1.3930 0.5020 ;
      RECT 1.0230 0.4100 1.3930 0.4600 ;
      RECT 1.3430 0.5020 1.7370 0.5520 ;
      RECT 1.6870 0.5520 1.7370 0.6780 ;
      RECT 1.6500 0.7280 1.7370 0.7520 ;
      RECT 1.6500 0.7520 1.7000 1.0200 ;
      RECT 1.0230 1.0200 1.7000 1.0700 ;
      RECT 3.3730 1.3900 5.5890 1.4400 ;
      RECT 3.9870 0.6670 4.3730 0.7170 ;
      RECT 2.1030 0.6130 2.5490 0.6630 ;
      RECT 2.1030 0.8670 2.8530 0.9170 ;
      RECT 2.1030 0.4130 2.1530 0.6130 ;
      RECT 2.1030 0.6630 2.1530 0.8670 ;
      RECT 5.2950 0.7310 5.3880 0.7810 ;
      RECT 5.2950 0.5050 5.3450 0.7310 ;
      RECT 5.3380 0.7810 5.3880 0.8670 ;
      RECT 5.3380 0.8670 5.5890 0.9170 ;
      RECT 5.3380 0.9170 5.3880 1.0320 ;
      RECT 5.2950 1.0320 5.3880 1.0820 ;
      RECT 5.2950 1.0820 5.3450 1.2400 ;
      RECT 8.2430 1.2000 9.3890 1.2500 ;
      RECT 0.7190 0.9410 0.9530 0.9910 ;
      RECT 3.8870 0.8670 4.1690 0.9170 ;
      RECT 4.1190 0.9170 4.1690 1.1270 ;
      RECT 3.0150 1.1270 4.1690 1.1770 ;
      RECT 3.0150 1.1770 3.0650 1.2400 ;
      RECT 3.0150 1.0660 3.1150 1.1270 ;
      RECT 3.0650 0.9170 3.1150 1.0660 ;
      RECT 3.0150 0.4130 3.0650 0.8670 ;
      RECT 3.0150 0.8670 3.3090 0.9170 ;
      RECT 3.8870 0.6070 3.9370 0.8670 ;
      RECT 3.8870 0.5570 3.9770 0.6070 ;
      RECT 3.9270 0.4130 3.9770 0.5570 ;
      RECT 2.5430 0.5130 2.6850 0.5630 ;
      RECT 2.6350 0.5630 2.6850 0.6130 ;
      RECT 2.6350 0.6130 2.8680 0.6630 ;
      RECT 2.6350 0.6630 2.6850 0.7540 ;
      RECT 2.5420 0.7540 2.6850 0.8040 ;
      RECT 1.1750 1.1330 1.5610 1.1830 ;
      RECT 0.7190 0.5100 1.2570 0.5600 ;
      RECT 0.8870 0.3100 1.5450 0.3600 ;
      RECT 1.4950 0.3600 1.5450 0.3920 ;
      RECT 0.8870 0.3600 0.9370 0.3920 ;
      RECT 3.4710 0.9670 4.0690 1.0170 ;
      RECT 3.1670 0.4070 3.2170 0.6190 ;
      RECT 3.4710 1.0170 3.5210 1.0770 ;
      RECT 3.4710 0.6690 3.5210 0.9670 ;
      RECT 3.1670 0.6190 3.5210 0.6690 ;
      RECT 3.4710 0.4070 3.5210 0.6190 ;
      RECT 4.5950 0.6130 4.8290 0.6630 ;
      RECT 2.6190 1.5240 4.8290 1.5740 ;
      RECT 2.3150 0.0940 4.5250 0.1440 ;
      RECT 4.4430 0.8670 4.6970 0.9170 ;
      RECT 7.0270 0.6130 7.3950 0.6630 ;
      RECT 7.3450 0.5700 7.3950 0.6130 ;
      RECT 7.3450 0.5200 7.8350 0.5700 ;
      RECT 7.7850 0.5700 7.8350 0.6040 ;
      RECT 7.7850 0.6040 8.0210 0.6540 ;
      RECT 8.7910 1.0620 9.2370 1.1120 ;
      RECT 8.7910 0.1260 8.8410 1.0620 ;
      RECT 1.4520 0.6020 1.6370 0.6520 ;
      RECT 0.2050 0.5260 0.2550 0.8410 ;
      RECT 0.2790 0.8910 0.3290 1.2140 ;
      RECT 0.2050 0.4760 0.3290 0.5260 ;
      RECT 0.2790 0.3160 0.3290 0.4760 ;
      RECT 0.2050 0.8410 1.5020 0.8910 ;
    LAYER PO ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 9.7890 0.0660 9.8190 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 8.2690 0.0670 8.2990 1.6050 ;
      RECT 3.7090 0.9390 3.7390 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
      RECT 3.7090 0.0660 3.7390 0.6370 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 2.7970 0.0660 2.8270 0.6910 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 11.0050 0.0660 11.0350 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 4.1650 0.9390 4.1950 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 10.8530 0.0660 10.8830 1.6060 ;
      RECT 9.4850 0.0660 9.5150 1.6060 ;
      RECT 5.9890 0.0660 6.0190 0.6910 ;
      RECT 10.7010 0.0660 10.7310 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 10.3970 0.0660 10.4270 1.6060 ;
      RECT 6.4450 0.0660 6.4750 0.7910 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 10.5490 0.0660 10.5790 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 10.0930 0.0660 10.1230 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 4.6210 0.0660 4.6510 0.6910 ;
      RECT 4.1650 0.0660 4.1950 0.6370 ;
      RECT 2.7970 0.8390 2.8270 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 6.4450 0.9390 6.4750 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 4.6210 0.8390 4.6510 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 9.3330 0.0660 9.3630 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6140 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 9.9410 0.0660 9.9710 1.6060 ;
      RECT 9.6370 0.0660 9.6670 1.6060 ;
      RECT 10.2450 0.0660 10.2750 1.6060 ;
      RECT 5.9890 0.9590 6.0190 1.6060 ;
    LAYER NWELL ;
      RECT -0.1160 1.5430 11.2040 1.7730 ;
      RECT -0.1160 0.6790 8.1620 1.5430 ;
      RECT 10.9290 0.6790 11.2040 1.5430 ;
      RECT 8.6230 0.4910 10.4690 1.0830 ;
  END
END RSDFFNARX2_LVT

MACRO RSDFFNSRARX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.032 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3770 1.4650 2.5490 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 10.0320 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 2.1030 1.1310 2.1530 1.6420 ;
        RECT 1.7990 1.1310 1.8490 1.6420 ;
        RECT 1.6470 1.1310 1.6970 1.6420 ;
        RECT 2.2550 1.2940 2.3050 1.6420 ;
        RECT 3.9670 1.2700 4.0170 1.6420 ;
        RECT 8.0710 1.4540 8.1210 1.6420 ;
        RECT 2.2550 1.2440 2.7770 1.2940 ;
        RECT 3.7580 1.2200 4.9050 1.2700 ;
        RECT 5.5990 1.4040 8.1210 1.4540 ;
        RECT 5.5990 1.2790 5.6490 1.4040 ;
        RECT 6.6630 0.9590 6.7130 1.4040 ;
        RECT 6.2070 0.9530 6.2570 1.4040 ;
    END
  END VDD

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.5110 0.4010 7.2110 0.4510 ;
        RECT 6.5110 0.1570 6.5610 0.4010 ;
        RECT 7.0890 0.4510 7.2110 0.5380 ;
        RECT 7.1610 0.5380 7.2110 0.8590 ;
        RECT 6.5110 0.8590 7.2110 0.9090 ;
        RECT 6.5110 0.9090 6.5610 1.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.8150 0.9690 7.3490 1.0190 ;
        RECT 7.2990 0.3510 7.3490 0.9690 ;
        RECT 6.8150 1.0190 7.0470 1.1290 ;
        RECT 6.7990 0.3010 7.3490 0.3510 ;
        RECT 6.8150 1.1290 6.8650 1.3270 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 10.0320 0.0300 ;
        RECT 2.1030 0.0300 2.1530 0.2970 ;
        RECT 9.0950 0.0300 9.1450 0.4260 ;
        RECT 1.6470 0.0300 1.6970 0.4050 ;
        RECT 6.6630 0.0300 6.7130 0.2410 ;
        RECT 1.7990 0.0300 1.8490 0.4050 ;
        RECT 7.7270 0.0300 7.7770 0.4260 ;
        RECT 0.5830 0.0300 0.6330 0.5120 ;
        RECT 0.4310 0.0300 0.4810 0.4340 ;
        RECT 8.6390 0.0300 8.6890 0.1980 ;
        RECT 6.3830 0.0300 6.4330 0.3000 ;
        RECT 2.1030 0.2970 3.9770 0.3470 ;
        RECT 5.5830 0.3000 6.4330 0.3500 ;
        RECT 3.7750 0.3470 3.8250 0.5570 ;
        RECT 2.5590 0.3470 2.6090 0.5570 ;
        RECT 2.7110 0.3470 2.7610 0.5570 ;
        RECT 2.1030 0.3470 2.1530 0.4050 ;
        RECT 3.9270 0.2380 3.9770 0.2970 ;
        RECT 3.9270 0.1880 4.9050 0.2380 ;
        RECT 4.2310 0.2380 4.2810 0.3490 ;
    END
  END VSS

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4390 0.0880 5.6890 0.1380 ;
        RECT 3.4390 0.1380 3.5970 0.2100 ;
        RECT 5.6390 0.1380 5.6890 0.2000 ;
        RECT 5.6390 0.2000 6.1810 0.2500 ;
        RECT 6.1310 0.0880 6.1810 0.2000 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.2170 0.2490 9.3290 0.3590 ;
        RECT 9.2280 0.3590 9.2780 0.5270 ;
        RECT 9.0030 0.5270 9.2780 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.5050 0.7050 4.6610 0.7310 ;
        RECT 4.5050 0.7310 4.9650 0.7810 ;
        RECT 4.6110 0.5970 4.6610 0.7050 ;
        RECT 4.5050 0.7810 4.6610 0.8150 ;
        RECT 4.9150 0.7810 4.9650 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 7.7110 0.9420 9.3290 1.0020 ;
        RECT 9.2190 0.6900 9.3290 0.9420 ;
        RECT 9.0950 0.6270 9.1450 0.9420 ;
    END
  END VDDG

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2520 1.3330 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6780 0.7250 0.7280 ;
        RECT 0.4010 0.5510 0.5110 0.6780 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 1.1610 1.0110 1.3160 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D
  OBS
    LAYER M1 ;
      RECT 5.1430 1.0170 5.1930 1.1200 ;
      RECT 5.1430 1.1700 5.1930 1.2700 ;
      RECT 4.6710 1.1200 5.1930 1.1700 ;
      RECT 4.1210 0.8580 4.2210 0.9080 ;
      RECT 4.1210 0.9080 4.1710 0.9680 ;
      RECT 3.6830 0.9680 4.1710 1.0180 ;
      RECT 1.4520 0.6020 1.6370 0.6520 ;
      RECT 0.2050 0.8410 1.5020 0.8910 ;
      RECT 1.4520 0.6520 1.5020 0.8410 ;
      RECT 0.2050 0.5260 0.2550 0.8410 ;
      RECT 0.2790 0.8910 0.3290 1.2140 ;
      RECT 0.2050 0.4760 0.3290 0.5260 ;
      RECT 0.2790 0.3160 0.3290 0.4760 ;
      RECT 3.1670 0.8540 4.0690 0.9040 ;
      RECT 3.1670 0.6130 3.2170 0.8540 ;
      RECT 3.1670 0.9040 3.2170 1.0590 ;
      RECT 3.1670 0.5630 3.3690 0.6130 ;
      RECT 3.1670 1.0590 3.5370 1.1090 ;
      RECT 3.3190 0.4070 3.3690 0.5630 ;
      RECT 3.1670 0.4130 3.2170 0.5630 ;
      RECT 3.1670 1.1090 3.2170 1.3370 ;
      RECT 6.2620 0.6320 6.6370 0.6820 ;
      RECT 6.5870 0.5970 6.6370 0.6320 ;
      RECT 5.8180 0.7290 6.0050 0.7790 ;
      RECT 5.9550 0.7790 6.0050 1.1790 ;
      RECT 5.8180 0.4500 5.8680 0.7290 ;
      RECT 5.4480 1.1790 6.0050 1.2290 ;
      RECT 6.2830 0.4500 6.3330 0.6320 ;
      RECT 5.4470 0.4000 6.3330 0.4500 ;
      RECT 5.4480 1.2290 5.4980 1.3530 ;
      RECT 5.4470 0.4500 5.4970 0.5630 ;
      RECT 5.4470 0.2970 5.4970 0.4000 ;
      RECT 2.9990 0.4120 3.1050 0.4620 ;
      RECT 3.0550 0.4620 3.1050 0.8130 ;
      RECT 3.0150 0.8130 3.1050 0.8630 ;
      RECT 3.0150 0.8630 3.0650 1.0830 ;
      RECT 2.2550 1.0830 3.0650 1.1330 ;
      RECT 3.0150 1.1330 3.0650 1.3540 ;
      RECT 2.2550 0.7520 2.3050 1.0830 ;
      RECT 2.2550 0.7020 2.3450 0.7520 ;
      RECT 2.2950 0.5510 2.3450 0.7020 ;
      RECT 2.2550 0.5010 2.3450 0.5510 ;
      RECT 2.2550 0.4070 2.3050 0.5010 ;
      RECT 2.4070 0.6130 2.8530 0.6630 ;
      RECT 2.4070 0.6630 2.4570 1.0040 ;
      RECT 2.4070 0.4130 2.4570 0.6130 ;
      RECT 8.0150 0.8200 8.5630 0.8700 ;
      RECT 1.6500 0.7020 1.9410 0.7280 ;
      RECT 1.6870 0.6780 1.9410 0.7020 ;
      RECT 1.3430 0.4600 1.3930 0.5020 ;
      RECT 1.0230 0.4100 1.3930 0.4600 ;
      RECT 1.0230 1.0200 1.7000 1.0700 ;
      RECT 1.6500 0.7520 1.7000 1.0200 ;
      RECT 1.6500 0.7280 1.7370 0.7520 ;
      RECT 1.6870 0.5520 1.7370 0.6780 ;
      RECT 1.3430 0.5020 1.7370 0.5520 ;
      RECT 0.8870 0.3100 1.5450 0.3600 ;
      RECT 1.4950 0.3600 1.5450 0.3920 ;
      RECT 0.8870 0.3600 0.9370 0.3920 ;
      RECT 5.5070 0.8660 5.6560 0.9160 ;
      RECT 5.6060 0.9160 5.6560 0.9670 ;
      RECT 5.6060 0.9670 5.7410 1.0170 ;
      RECT 6.6870 0.6130 7.1090 0.6630 ;
      RECT 6.0550 0.8090 6.1050 1.3010 ;
      RECT 6.0550 0.6780 6.1050 0.7590 ;
      RECT 5.9630 0.6280 6.1050 0.6780 ;
      RECT 6.0550 0.5000 6.1050 0.6280 ;
      RECT 6.3590 0.8090 6.4090 1.3010 ;
      RECT 6.6870 0.6630 6.7370 0.7590 ;
      RECT 6.0550 0.7590 6.7370 0.8090 ;
      RECT 1.9910 0.6280 2.2450 0.6520 ;
      RECT 1.9520 0.6020 2.2450 0.6280 ;
      RECT 1.9910 0.6520 2.0410 0.7780 ;
      RECT 1.9520 0.5780 2.0410 0.6020 ;
      RECT 1.9520 0.7780 2.0410 0.8280 ;
      RECT 1.9520 0.3190 2.0020 0.5780 ;
      RECT 1.9520 0.8280 2.0020 1.0760 ;
      RECT 8.3190 0.7090 8.8570 0.7590 ;
      RECT 5.0310 0.5380 5.0810 1.0200 ;
      RECT 4.5190 0.5110 5.0810 0.5380 ;
      RECT 4.5350 1.0200 5.0810 1.0700 ;
      RECT 4.5190 0.4880 5.0800 0.5110 ;
      RECT 4.2710 0.7880 4.3210 1.1200 ;
      RECT 3.3740 0.7380 4.3230 0.7880 ;
      RECT 4.0790 0.5050 4.1290 0.7380 ;
      RECT 4.5350 1.0700 4.5850 1.1200 ;
      RECT 4.0580 1.1200 4.5850 1.1700 ;
      RECT 8.9430 0.6770 8.9930 0.7680 ;
      RECT 8.9030 0.4270 8.9930 0.4620 ;
      RECT 8.9430 0.1260 8.9930 0.4270 ;
      RECT 8.9030 0.6270 8.9930 0.6770 ;
      RECT 8.9030 0.5120 8.9530 0.6270 ;
      RECT 8.6990 0.4770 8.9530 0.5120 ;
      RECT 8.6990 0.4620 8.9930 0.4770 ;
      RECT 2.9220 0.0940 3.3150 0.1440 ;
      RECT 4.2910 1.5200 4.9810 1.5700 ;
      RECT 4.7460 0.6130 4.9810 0.6630 ;
      RECT 5.2950 0.8670 5.4370 0.9170 ;
      RECT 5.2950 0.6630 5.3450 0.8670 ;
      RECT 5.2950 0.6130 5.7410 0.6630 ;
      RECT 4.3830 0.9200 4.8130 0.9700 ;
      RECT 4.7630 0.8310 4.8130 0.9200 ;
      RECT 4.3830 0.9700 4.4330 1.0340 ;
      RECT 4.3830 0.5050 4.4330 0.9200 ;
      RECT 4.1390 1.4200 5.4450 1.4700 ;
      RECT 3.3030 1.1900 3.6890 1.2400 ;
      RECT 3.2270 1.3890 3.7650 1.4390 ;
      RECT 4.9950 0.1880 5.5890 0.2380 ;
      RECT 4.9950 0.2380 5.0450 0.2880 ;
      RECT 4.3540 0.2880 5.0450 0.3380 ;
      RECT 3.9470 0.4550 3.9970 0.6130 ;
      RECT 3.6830 0.6130 3.9970 0.6630 ;
      RECT 4.3540 0.3380 4.4040 0.4050 ;
      RECT 3.9470 0.4050 4.4040 0.4550 ;
      RECT 7.0270 1.1990 8.3250 1.2490 ;
      RECT 2.6190 1.5240 3.9170 1.5740 ;
      RECT 8.3190 0.1320 8.5530 0.1820 ;
      RECT 7.5750 1.0620 8.0240 1.1120 ;
      RECT 7.5750 0.6770 7.6250 1.0620 ;
      RECT 7.5350 0.6270 7.6250 0.6770 ;
      RECT 7.5350 0.4770 7.5850 0.6270 ;
      RECT 7.5350 0.4270 7.6250 0.4770 ;
      RECT 7.5750 0.1260 7.6250 0.4270 ;
      RECT 7.6350 0.5270 8.2330 0.5770 ;
      RECT 7.8790 0.5770 7.9290 0.8840 ;
      RECT 7.8790 0.1260 7.9290 0.5270 ;
      RECT 8.1830 0.5770 8.2330 0.7700 ;
      RECT 8.1830 0.3480 8.2330 0.5270 ;
      RECT 5.8110 0.0940 6.0450 0.1440 ;
      RECT 0.7190 0.5100 1.2570 0.5600 ;
      RECT 1.1750 1.1330 1.5610 1.1830 ;
      RECT 0.7190 0.9410 0.9530 0.9910 ;
      RECT 8.5470 1.0620 9.0850 1.1120 ;
      RECT 8.0150 0.2480 8.8570 0.2980 ;
      RECT 5.0490 1.5200 8.0210 1.5700 ;
      RECT 2.8630 0.7130 2.9890 0.7630 ;
      RECT 2.8630 0.7630 2.9130 1.0330 ;
      RECT 2.9390 0.5630 2.9890 0.7130 ;
      RECT 2.8470 0.5130 2.9890 0.5630 ;
      RECT 4.6710 0.3880 5.3450 0.4380 ;
      RECT 5.2950 0.4380 5.3450 0.5630 ;
      RECT 5.2950 0.2970 5.3450 0.3880 ;
      RECT 5.1430 0.4380 5.1930 0.9670 ;
      RECT 5.1430 0.9670 5.3610 1.0170 ;
    LAYER PO ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 5.6850 0.0660 5.7150 0.6910 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 3.1010 0.8400 3.1310 1.6060 ;
      RECT 5.6850 0.9390 5.7150 1.6060 ;
      RECT 5.3810 0.0660 5.4110 0.6370 ;
      RECT 3.1010 0.0660 3.1310 0.6370 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 3.7090 0.0660 3.7390 0.6910 ;
      RECT 4.9250 0.0660 4.9550 0.6910 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 9.3330 0.0660 9.3630 1.6060 ;
      RECT 4.6210 0.8920 4.6510 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 5.3810 0.8390 5.4110 1.6060 ;
      RECT 9.4850 0.0660 9.5150 1.6060 ;
      RECT 9.9410 0.0660 9.9710 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 9.6370 0.0660 9.6670 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 9.7890 0.0660 9.8190 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 4.6210 0.0660 4.6510 0.6910 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 3.7090 0.9390 3.7390 1.6060 ;
      RECT 7.0530 0.0670 7.0830 1.6050 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 4.9250 0.8390 4.9550 1.6060 ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
    LAYER NWELL ;
      RECT 7.4080 0.4910 9.4190 1.0830 ;
      RECT -0.1150 1.5430 10.1540 1.7730 ;
      RECT -0.1150 0.6790 6.9460 1.5430 ;
      RECT 9.8790 0.6790 10.1540 1.5430 ;
  END
END RSDFFNSRARX1_LVT

MACRO RSDFFNSRARX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.336 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3770 1.4650 2.5490 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 10.3360 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 2.1030 1.1310 2.1530 1.6420 ;
        RECT 1.7990 1.1310 1.8490 1.6420 ;
        RECT 1.6470 1.1310 1.6970 1.6420 ;
        RECT 8.3750 1.4540 8.4250 1.6420 ;
        RECT 2.2550 1.2940 2.3050 1.6420 ;
        RECT 3.9670 1.2700 4.0170 1.6420 ;
        RECT 5.5990 1.4040 8.4250 1.4540 ;
        RECT 2.2550 1.2440 2.7770 1.2940 ;
        RECT 3.7580 1.2200 4.9050 1.2700 ;
        RECT 5.5990 1.2790 5.6490 1.4040 ;
        RECT 6.2070 0.9530 6.2570 1.4040 ;
        RECT 6.8150 0.9610 6.8650 1.4040 ;
        RECT 7.1190 1.0530 7.1690 1.4040 ;
        RECT 6.5110 0.9130 6.5610 1.4040 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 10.3360 0.0300 ;
        RECT 2.1030 0.0300 2.1530 0.2970 ;
        RECT 6.8150 0.0300 6.8650 0.3200 ;
        RECT 9.3990 0.0300 9.4490 0.4260 ;
        RECT 1.6470 0.0300 1.6970 0.4050 ;
        RECT 6.5110 0.0300 6.5610 0.4090 ;
        RECT 7.1190 0.0300 7.1690 0.2210 ;
        RECT 1.7990 0.0300 1.8490 0.4050 ;
        RECT 8.0310 0.0300 8.0810 0.4260 ;
        RECT 0.5830 0.0300 0.6330 0.5120 ;
        RECT 0.4310 0.0300 0.4810 0.4340 ;
        RECT 8.9430 0.0300 8.9930 0.1980 ;
        RECT 6.3830 0.0300 6.4330 0.3000 ;
        RECT 2.1030 0.2970 3.9770 0.3470 ;
        RECT 5.5830 0.3000 6.4330 0.3500 ;
        RECT 3.7750 0.3470 3.8250 0.5570 ;
        RECT 2.5590 0.3470 2.6090 0.5570 ;
        RECT 2.7110 0.3470 2.7610 0.5570 ;
        RECT 2.1030 0.3470 2.1530 0.4050 ;
        RECT 3.9270 0.2380 3.9770 0.2970 ;
        RECT 3.9270 0.1880 4.9050 0.2380 ;
        RECT 4.2310 0.2380 4.2810 0.3490 ;
    END
  END VSS

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4390 0.0880 5.6890 0.1380 ;
        RECT 3.4390 0.1380 3.5970 0.2100 ;
        RECT 5.6390 0.1380 5.6890 0.2000 ;
        RECT 5.6390 0.2000 6.1810 0.2500 ;
        RECT 6.1310 0.0880 6.1810 0.2000 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.5210 0.2490 9.6310 0.3590 ;
        RECT 9.5320 0.3590 9.5820 0.5270 ;
        RECT 9.3070 0.5270 9.5820 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.5050 0.7160 4.6610 0.7310 ;
        RECT 4.5050 0.7310 4.9650 0.7810 ;
        RECT 4.6110 0.5970 4.6610 0.7160 ;
        RECT 4.5050 0.7810 4.6610 0.8150 ;
        RECT 4.9150 0.7810 4.9650 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.6630 0.1490 6.7130 0.4020 ;
        RECT 6.6630 0.4020 7.5150 0.4520 ;
        RECT 7.3930 0.4520 7.5150 0.5120 ;
        RECT 7.4650 0.5120 7.5150 0.8330 ;
        RECT 6.6630 0.8330 7.5150 0.8830 ;
        RECT 6.6630 0.8830 6.7130 1.3190 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.9670 0.2710 7.6650 0.3210 ;
        RECT 7.5450 0.3210 7.6650 0.3600 ;
        RECT 7.5450 0.2500 7.6650 0.2710 ;
        RECT 6.9670 0.1490 7.0170 0.2710 ;
        RECT 7.6150 0.3600 7.6650 0.9330 ;
        RECT 7.5450 0.2490 7.6550 0.2500 ;
        RECT 6.9670 0.9330 7.6650 0.9830 ;
        RECT 6.9670 0.9830 7.0170 1.3270 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 8.0150 0.9420 9.6330 1.0020 ;
        RECT 9.5230 0.6900 9.6330 0.9420 ;
        RECT 9.3990 0.6270 9.4490 0.9420 ;
    END
  END VDDG

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2520 1.3330 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6780 0.7250 0.7280 ;
        RECT 0.4010 0.5510 0.5110 0.6780 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 1.1610 1.0110 1.3160 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D
  OBS
    LAYER M1 ;
      RECT 5.1430 1.1700 5.1930 1.2700 ;
      RECT 4.6710 1.1200 5.1930 1.1700 ;
      RECT 4.1210 0.8580 4.2210 0.9080 ;
      RECT 4.1210 0.9080 4.1710 0.9680 ;
      RECT 3.6830 0.9680 4.1710 1.0180 ;
      RECT 1.4520 0.6020 1.6370 0.6520 ;
      RECT 0.2050 0.8410 1.5020 0.8910 ;
      RECT 1.4520 0.6520 1.5020 0.8410 ;
      RECT 0.2050 0.5260 0.2550 0.8410 ;
      RECT 0.2790 0.8910 0.3290 1.2140 ;
      RECT 0.2050 0.4760 0.3290 0.5260 ;
      RECT 0.2790 0.3160 0.3290 0.4760 ;
      RECT 6.8680 0.6130 7.4130 0.6630 ;
      RECT 6.8680 0.6630 6.9180 0.7320 ;
      RECT 6.0550 0.7320 6.9180 0.7820 ;
      RECT 6.0550 0.7820 6.1050 1.3010 ;
      RECT 6.0550 0.6780 6.1050 0.7320 ;
      RECT 5.9630 0.6280 6.1050 0.6780 ;
      RECT 6.0550 0.5000 6.1050 0.6280 ;
      RECT 6.3590 0.7820 6.4090 1.3010 ;
      RECT 3.1670 0.8540 4.0690 0.9040 ;
      RECT 3.3190 0.4070 3.3690 0.5630 ;
      RECT 3.1670 0.5630 3.3690 0.6130 ;
      RECT 3.1670 0.4130 3.2170 0.5630 ;
      RECT 3.1670 0.6130 3.2170 0.8540 ;
      RECT 3.1670 0.9040 3.2170 1.0590 ;
      RECT 3.1670 1.0590 3.5370 1.1090 ;
      RECT 3.1670 1.1090 3.2170 1.3370 ;
      RECT 6.2620 0.6320 6.8050 0.6820 ;
      RECT 5.8180 0.4500 5.8680 0.7290 ;
      RECT 5.8180 0.7290 6.0050 0.7790 ;
      RECT 5.9550 0.7790 6.0050 1.1790 ;
      RECT 5.4480 1.1790 6.0050 1.2290 ;
      RECT 6.2830 0.4500 6.3330 0.6320 ;
      RECT 5.4470 0.4000 6.3330 0.4500 ;
      RECT 5.4470 0.4500 5.4970 0.5630 ;
      RECT 5.4470 0.2970 5.4970 0.4000 ;
      RECT 5.4480 1.2290 5.4980 1.3530 ;
      RECT 4.9950 0.1880 5.5890 0.2380 ;
      RECT 4.9950 0.2380 5.0450 0.2880 ;
      RECT 4.3540 0.2880 5.0450 0.3380 ;
      RECT 3.9470 0.4550 3.9970 0.6130 ;
      RECT 3.6830 0.6130 3.9970 0.6630 ;
      RECT 4.3540 0.3380 4.4040 0.4050 ;
      RECT 3.9470 0.4050 4.4040 0.4550 ;
      RECT 3.0150 0.8130 3.1050 0.8630 ;
      RECT 3.0550 0.4620 3.1050 0.8130 ;
      RECT 3.0150 0.8630 3.0650 1.0830 ;
      RECT 2.9990 0.4120 3.1050 0.4620 ;
      RECT 2.2550 1.0830 3.0650 1.1330 ;
      RECT 3.0150 1.1330 3.0650 1.3540 ;
      RECT 2.2550 0.7520 2.3050 1.0830 ;
      RECT 2.2550 0.7020 2.3450 0.7520 ;
      RECT 2.2950 0.5510 2.3450 0.7020 ;
      RECT 2.2550 0.5010 2.3450 0.5510 ;
      RECT 2.2550 0.4070 2.3050 0.5010 ;
      RECT 2.4070 0.6130 2.8530 0.6630 ;
      RECT 2.4070 0.6630 2.4570 1.0040 ;
      RECT 2.4070 0.4130 2.4570 0.6130 ;
      RECT 8.3190 0.8200 8.8670 0.8700 ;
      RECT 1.6500 0.7020 1.9410 0.7280 ;
      RECT 1.6870 0.6780 1.9410 0.7020 ;
      RECT 1.3430 0.4600 1.3930 0.5020 ;
      RECT 1.0230 0.4100 1.3930 0.4600 ;
      RECT 1.0230 1.0200 1.7000 1.0700 ;
      RECT 1.6500 0.7520 1.7000 1.0200 ;
      RECT 1.6500 0.7280 1.7370 0.7520 ;
      RECT 1.6870 0.5520 1.7370 0.6780 ;
      RECT 1.3430 0.5020 1.7370 0.5520 ;
      RECT 0.8870 0.3100 1.5450 0.3600 ;
      RECT 1.4950 0.3600 1.5450 0.3920 ;
      RECT 0.8870 0.3600 0.9370 0.3920 ;
      RECT 5.5070 0.8660 5.6560 0.9160 ;
      RECT 5.6060 0.9160 5.6560 0.9670 ;
      RECT 5.6060 0.9670 5.7410 1.0170 ;
      RECT 1.9910 0.6280 2.2450 0.6520 ;
      RECT 1.9520 0.6020 2.2450 0.6280 ;
      RECT 1.9910 0.6520 2.0410 0.7780 ;
      RECT 1.9520 0.5780 2.0410 0.6020 ;
      RECT 1.9520 0.7780 2.0410 0.8280 ;
      RECT 1.9520 0.3190 2.0020 0.5780 ;
      RECT 1.9520 0.8280 2.0020 1.0760 ;
      RECT 8.6230 0.7090 9.1610 0.7590 ;
      RECT 8.8510 1.0620 9.3890 1.1120 ;
      RECT 8.3190 0.2480 9.1610 0.2980 ;
      RECT 5.0310 0.5380 5.0810 1.0200 ;
      RECT 4.5190 0.5110 5.0810 0.5380 ;
      RECT 4.5350 1.0200 5.0810 1.0700 ;
      RECT 4.5190 0.4880 5.0800 0.5110 ;
      RECT 4.2710 0.7880 4.3210 1.1200 ;
      RECT 3.3740 0.7380 4.3230 0.7880 ;
      RECT 4.0790 0.5050 4.1290 0.7380 ;
      RECT 4.5350 1.0700 4.5850 1.1200 ;
      RECT 4.0580 1.1200 4.5850 1.1700 ;
      RECT 5.0490 1.5200 8.3250 1.5700 ;
      RECT 9.2470 0.6770 9.2970 0.7680 ;
      RECT 9.2070 0.4270 9.2970 0.4620 ;
      RECT 9.2470 0.1260 9.2970 0.4270 ;
      RECT 9.2070 0.6270 9.2970 0.6770 ;
      RECT 9.2070 0.5120 9.2570 0.6270 ;
      RECT 9.0030 0.4770 9.2570 0.5120 ;
      RECT 9.0030 0.4620 9.2970 0.4770 ;
      RECT 2.9220 0.0940 3.3150 0.1440 ;
      RECT 4.2910 1.5200 4.9810 1.5700 ;
      RECT 4.7460 0.6130 4.9810 0.6630 ;
      RECT 5.2950 0.8670 5.4370 0.9170 ;
      RECT 5.2950 0.6630 5.3450 0.8670 ;
      RECT 5.2950 0.6130 5.7410 0.6630 ;
      RECT 4.3830 0.9200 4.8130 0.9700 ;
      RECT 4.7630 0.8310 4.8130 0.9200 ;
      RECT 4.3830 0.9700 4.4330 1.0340 ;
      RECT 4.3830 0.5050 4.4330 0.9200 ;
      RECT 4.1390 1.4200 5.4450 1.4700 ;
      RECT 3.3030 1.1900 3.6890 1.2400 ;
      RECT 3.2270 1.3890 3.7650 1.4390 ;
      RECT 7.3310 1.1990 8.6290 1.2490 ;
      RECT 7.9390 0.5270 8.5370 0.5770 ;
      RECT 8.4870 0.5770 8.5370 0.7700 ;
      RECT 8.4870 0.3480 8.5370 0.5270 ;
      RECT 8.1830 0.5770 8.2330 0.8800 ;
      RECT 8.1830 0.1260 8.2330 0.5270 ;
      RECT 2.6190 1.5240 3.9170 1.5740 ;
      RECT 8.6230 0.1320 8.8570 0.1820 ;
      RECT 7.8790 1.0630 8.3280 1.1130 ;
      RECT 7.8790 0.6770 7.9290 1.0630 ;
      RECT 7.8390 0.6270 7.9290 0.6770 ;
      RECT 7.8390 0.4770 7.8890 0.6270 ;
      RECT 7.8390 0.4270 7.9290 0.4770 ;
      RECT 7.8790 0.1260 7.9290 0.4270 ;
      RECT 5.8110 0.0940 6.0450 0.1440 ;
      RECT 0.7190 0.5100 1.2570 0.5600 ;
      RECT 1.1750 1.1330 1.5610 1.1830 ;
      RECT 0.7190 0.9410 0.9530 0.9910 ;
      RECT 2.8630 0.7130 2.9890 0.7630 ;
      RECT 2.8630 0.7630 2.9130 1.0330 ;
      RECT 2.9390 0.5630 2.9890 0.7130 ;
      RECT 2.8470 0.5130 2.9890 0.5630 ;
      RECT 4.6710 0.3880 5.3450 0.4380 ;
      RECT 5.2950 0.4380 5.3450 0.5630 ;
      RECT 5.2950 0.2970 5.3450 0.3880 ;
      RECT 5.1430 0.4380 5.1930 0.9670 ;
      RECT 5.1430 0.9670 5.3610 1.0170 ;
      RECT 5.1430 1.0170 5.1930 1.1200 ;
    LAYER PO ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 4.9250 0.8390 4.9550 1.6060 ;
      RECT 9.4850 0.0660 9.5150 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 5.6850 0.0660 5.7150 0.6910 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 3.1010 0.8400 3.1310 1.6060 ;
      RECT 5.6850 0.9390 5.7150 1.6060 ;
      RECT 5.3810 0.0660 5.4110 0.6370 ;
      RECT 3.1010 0.0660 3.1310 0.6370 ;
      RECT 9.3330 0.0660 9.3630 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 3.7090 0.0660 3.7390 0.6910 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 4.9250 0.0660 4.9550 0.6910 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 9.6370 0.0660 9.6670 1.6060 ;
      RECT 4.6210 0.8920 4.6510 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 5.3810 0.8390 5.4110 1.6060 ;
      RECT 9.7890 0.0660 9.8190 1.6060 ;
      RECT 10.2450 0.0660 10.2750 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 9.9410 0.0660 9.9710 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 10.0930 0.0660 10.1230 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 4.6210 0.0660 4.6510 0.6910 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 3.7090 0.9390 3.7390 1.6060 ;
      RECT 7.3570 0.0670 7.3870 1.6050 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
    LAYER NWELL ;
      RECT 7.7120 0.4910 9.7230 1.0830 ;
      RECT -0.1150 1.5430 10.4580 1.7730 ;
      RECT -0.1150 0.6790 7.2500 1.5430 ;
      RECT 10.1830 0.6790 10.4580 1.5430 ;
  END
END RSDFFNSRARX2_LVT

MACRO RSDFFNSRASRNX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.488 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 10.4880 1.7020 ;
        RECT 0.5830 1.0330 0.6330 1.6420 ;
        RECT 0.4310 1.0330 0.4810 1.6420 ;
        RECT 2.1030 1.1310 2.1530 1.6420 ;
        RECT 1.7990 1.1310 1.8490 1.6420 ;
        RECT 1.6470 1.1310 1.6970 1.6420 ;
        RECT 8.3750 1.4540 8.4250 1.6420 ;
        RECT 3.9670 1.2700 4.0170 1.6420 ;
        RECT 2.2550 1.2940 2.3050 1.6420 ;
        RECT 5.7510 1.4040 8.4250 1.4540 ;
        RECT 3.7580 1.2200 5.0570 1.2700 ;
        RECT 2.2550 1.2440 2.7770 1.2940 ;
        RECT 5.7510 1.2790 5.8010 1.4040 ;
        RECT 6.9670 0.9590 7.0170 1.4040 ;
        RECT 6.5110 0.9530 6.5610 1.4040 ;
    END
  END VDD

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.8150 0.4010 7.5150 0.4510 ;
        RECT 6.8150 0.1570 6.8650 0.4010 ;
        RECT 7.3930 0.4510 7.5150 0.5380 ;
        RECT 7.4650 0.5380 7.5150 0.8590 ;
        RECT 6.8150 0.8590 7.5150 0.9090 ;
        RECT 6.8150 0.9090 6.8650 1.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 10.4880 0.0300 ;
        RECT 2.1030 0.0300 2.1530 0.3070 ;
        RECT 9.3990 0.0300 9.4490 0.4260 ;
        RECT 1.6470 0.0300 1.6970 0.4050 ;
        RECT 6.9670 0.0300 7.0170 0.2410 ;
        RECT 1.7990 0.0300 1.8490 0.4050 ;
        RECT 8.0310 0.0300 8.0810 0.4260 ;
        RECT 0.5830 0.0300 0.6330 0.5120 ;
        RECT 0.4310 0.0300 0.4810 0.4340 ;
        RECT 8.9430 0.0300 8.9930 0.1980 ;
        RECT 6.6870 0.0300 6.7370 0.2880 ;
        RECT 2.1030 0.3070 3.9770 0.3570 ;
        RECT 5.7350 0.2880 6.7370 0.3380 ;
        RECT 2.5590 0.3570 2.6090 0.5570 ;
        RECT 3.7750 0.3570 3.8250 0.5570 ;
        RECT 2.7110 0.3570 2.7610 0.5570 ;
        RECT 3.9270 0.3570 3.9770 0.5330 ;
        RECT 2.1030 0.3570 2.1530 0.4050 ;
        RECT 3.9270 0.2380 3.9770 0.3070 ;
        RECT 3.9270 0.1880 5.0570 0.2380 ;
        RECT 4.3830 0.2380 4.4330 0.3490 ;
    END
  END VSS

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.9790 0.8570 6.1350 0.9750 ;
        RECT 5.9790 0.9750 6.0290 1.0790 ;
        RECT 5.4470 1.0790 6.0290 1.1290 ;
        RECT 5.4470 1.1290 5.4970 1.3200 ;
        RECT 4.1550 1.3200 5.4970 1.3700 ;
        RECT 4.1550 1.3700 4.2050 1.4550 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4390 0.0880 6.4850 0.1380 ;
        RECT 3.4390 0.1380 3.6370 0.2100 ;
        RECT 6.4350 0.1380 6.4850 0.1700 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3770 1.4650 2.5490 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.5210 0.2490 9.6310 0.3590 ;
        RECT 9.5320 0.3590 9.5820 0.5270 ;
        RECT 9.3070 0.5270 9.5820 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6570 0.7050 4.8130 0.7310 ;
        RECT 4.6570 0.7310 5.1170 0.7810 ;
        RECT 4.7630 0.5970 4.8130 0.7050 ;
        RECT 4.6570 0.7810 4.8130 0.8150 ;
        RECT 5.0670 0.7810 5.1170 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 8.0150 0.9490 9.6330 1.0090 ;
        RECT 9.5230 0.6900 9.6330 0.9490 ;
        RECT 9.3990 1.0090 9.4490 1.0170 ;
        RECT 9.3990 0.6270 9.4490 0.9490 ;
    END
  END VDDG

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2520 1.3330 1.4230 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SI

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6780 0.7250 0.7280 ;
        RECT 0.4010 0.5510 0.5110 0.6780 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 1.1610 1.0110 1.3160 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D
  OBS
    LAYER M1 ;
      RECT 5.2950 0.4380 5.3450 0.9670 ;
      RECT 5.2950 1.0170 5.3450 1.1200 ;
      RECT 5.2950 1.1700 5.3450 1.2700 ;
      RECT 4.8230 1.1200 5.3450 1.1700 ;
      RECT 4.2130 0.8580 4.3730 0.9080 ;
      RECT 4.2130 0.9080 4.2630 0.9680 ;
      RECT 3.6830 0.9680 4.2630 1.0180 ;
      RECT 1.4520 0.6020 1.6370 0.6520 ;
      RECT 0.2050 0.8410 1.5020 0.8910 ;
      RECT 1.4520 0.6520 1.5020 0.8410 ;
      RECT 0.2050 0.5260 0.2550 0.8410 ;
      RECT 0.2790 0.8910 0.3290 1.2140 ;
      RECT 0.2050 0.4760 0.3290 0.5260 ;
      RECT 0.2790 0.3160 0.3290 0.4760 ;
      RECT 3.1670 0.8540 4.0690 0.9040 ;
      RECT 3.1670 0.6130 3.2170 0.8540 ;
      RECT 3.1670 0.9040 3.2170 1.0590 ;
      RECT 3.1670 0.5630 3.3690 0.6130 ;
      RECT 3.1670 1.0590 3.5370 1.1090 ;
      RECT 3.3190 0.4070 3.3690 0.5630 ;
      RECT 3.1670 0.4130 3.2170 0.5630 ;
      RECT 3.1670 1.1090 3.2170 1.3370 ;
      RECT 6.5870 0.6420 6.9410 0.6920 ;
      RECT 6.8910 0.5970 6.9410 0.6420 ;
      RECT 5.9430 0.7290 6.3090 0.7790 ;
      RECT 6.2590 0.7790 6.3090 1.1790 ;
      RECT 5.9430 0.4500 5.9930 0.7290 ;
      RECT 5.5990 0.4000 6.6370 0.4500 ;
      RECT 6.5870 0.4500 6.6370 0.6420 ;
      RECT 5.6000 1.1790 6.3090 1.2290 ;
      RECT 5.6000 1.2290 5.6500 1.3530 ;
      RECT 5.5990 0.4500 5.6490 0.5630 ;
      RECT 5.5990 0.2970 5.6490 0.4000 ;
      RECT 3.0150 0.8130 3.1050 0.8630 ;
      RECT 3.0550 0.4620 3.1050 0.8130 ;
      RECT 3.0150 0.8630 3.0650 1.0830 ;
      RECT 2.9990 0.4120 3.1050 0.4620 ;
      RECT 2.2550 1.0830 3.0650 1.1330 ;
      RECT 3.0150 1.1330 3.0650 1.3540 ;
      RECT 2.2550 0.7520 2.3050 1.0830 ;
      RECT 2.2550 0.7020 2.3450 0.7520 ;
      RECT 2.2950 0.5510 2.3450 0.7020 ;
      RECT 2.2550 0.5010 2.3450 0.5510 ;
      RECT 2.2550 0.4070 2.3050 0.5010 ;
      RECT 2.4070 0.6130 2.8530 0.6630 ;
      RECT 2.4070 0.6630 2.4570 1.0040 ;
      RECT 2.4070 0.4130 2.4570 0.6130 ;
      RECT 8.3190 0.8200 8.8670 0.8700 ;
      RECT 1.6500 0.7020 1.9410 0.7280 ;
      RECT 1.6870 0.6780 1.9410 0.7020 ;
      RECT 1.3430 0.4600 1.3930 0.5020 ;
      RECT 1.0230 0.4100 1.3930 0.4600 ;
      RECT 1.0230 1.0200 1.7000 1.0700 ;
      RECT 1.6500 0.7520 1.7000 1.0200 ;
      RECT 1.6500 0.7280 1.7370 0.7520 ;
      RECT 1.6870 0.5520 1.7370 0.6780 ;
      RECT 1.3430 0.5020 1.7370 0.5520 ;
      RECT 0.8870 0.3100 1.5450 0.3600 ;
      RECT 1.4950 0.3600 1.5450 0.3920 ;
      RECT 0.8870 0.3600 0.9370 0.3920 ;
      RECT 5.6590 0.8660 5.8080 0.9160 ;
      RECT 5.7580 0.9160 5.8080 0.9670 ;
      RECT 5.7580 0.9670 5.8930 1.0170 ;
      RECT 6.9910 0.6130 7.4130 0.6630 ;
      RECT 6.3590 0.8090 6.4090 1.3010 ;
      RECT 6.3590 0.5500 6.4090 0.7590 ;
      RECT 6.1310 0.5000 6.4090 0.5500 ;
      RECT 6.1310 0.5500 6.1810 0.6790 ;
      RECT 6.6630 0.8090 6.7130 1.3010 ;
      RECT 6.9910 0.6630 7.0410 0.7590 ;
      RECT 6.3590 0.7590 7.0410 0.8090 ;
      RECT 1.9910 0.6280 2.2450 0.6520 ;
      RECT 1.9520 0.6020 2.2450 0.6280 ;
      RECT 1.9910 0.6520 2.0410 0.7780 ;
      RECT 1.9520 0.5780 2.0410 0.6020 ;
      RECT 1.9520 0.7780 2.0410 0.8280 ;
      RECT 1.9520 0.3190 2.0020 0.5780 ;
      RECT 1.9520 0.8280 2.0020 1.0760 ;
      RECT 8.6230 0.7090 9.1610 0.7590 ;
      RECT 5.2010 1.5200 8.3250 1.5700 ;
      RECT 5.1830 0.5380 5.2330 1.0200 ;
      RECT 4.6710 0.5070 5.2330 0.5380 ;
      RECT 4.6870 1.0200 5.2330 1.0700 ;
      RECT 4.6710 0.4880 5.2320 0.5070 ;
      RECT 4.4230 0.7880 4.4730 1.1200 ;
      RECT 3.3740 0.7380 4.4750 0.7880 ;
      RECT 4.2310 0.5050 4.2810 0.7380 ;
      RECT 4.6870 1.0700 4.7370 1.1200 ;
      RECT 3.9110 1.1200 4.7370 1.1700 ;
      RECT 9.2470 0.6770 9.2970 0.7680 ;
      RECT 9.2070 0.4270 9.2970 0.4620 ;
      RECT 9.2470 0.1260 9.2970 0.4270 ;
      RECT 9.2070 0.6270 9.2970 0.6770 ;
      RECT 9.2070 0.5120 9.2570 0.6270 ;
      RECT 9.0030 0.4770 9.2570 0.5120 ;
      RECT 9.0030 0.4620 9.2970 0.4770 ;
      RECT 2.9220 0.0940 3.3150 0.1440 ;
      RECT 4.4430 1.5200 5.1330 1.5700 ;
      RECT 4.8980 0.6130 5.1330 0.6630 ;
      RECT 5.4470 0.8670 5.5890 0.9170 ;
      RECT 5.4470 0.6630 5.4970 0.8670 ;
      RECT 5.4470 0.6130 5.8930 0.6630 ;
      RECT 4.5350 0.9200 4.9650 0.9700 ;
      RECT 4.9150 0.8310 4.9650 0.9200 ;
      RECT 4.5350 0.9700 4.5850 1.0340 ;
      RECT 4.5350 0.5050 4.5850 0.9200 ;
      RECT 4.2910 1.4200 5.5970 1.4700 ;
      RECT 3.3030 1.1900 3.6890 1.2400 ;
      RECT 5.8800 1.2870 6.2730 1.3370 ;
      RECT 3.2270 1.3890 3.7650 1.4390 ;
      RECT 5.1470 0.1880 5.7410 0.2380 ;
      RECT 5.1470 0.2380 5.1970 0.2880 ;
      RECT 4.5060 0.2880 5.1970 0.3380 ;
      RECT 4.1190 0.4550 4.1690 0.6130 ;
      RECT 3.6830 0.6130 4.1690 0.6630 ;
      RECT 4.5060 0.3380 4.5560 0.4050 ;
      RECT 4.1190 0.4050 4.5560 0.4550 ;
      RECT 2.6190 1.5240 3.9170 1.5740 ;
      RECT 7.3310 1.2690 8.6290 1.3190 ;
      RECT 7.9390 0.5270 8.5370 0.5770 ;
      RECT 8.4870 0.5770 8.5370 0.7700 ;
      RECT 8.4870 0.3480 8.5370 0.5270 ;
      RECT 8.1830 0.5770 8.2330 0.8790 ;
      RECT 8.1830 0.1260 8.2330 0.5270 ;
      RECT 8.6230 0.1320 8.8570 0.1820 ;
      RECT 7.8790 1.1370 8.3280 1.1870 ;
      RECT 7.8790 0.6770 7.9290 1.1370 ;
      RECT 7.8390 0.6270 7.9290 0.6770 ;
      RECT 7.8390 0.4770 7.8890 0.6270 ;
      RECT 7.8390 0.4270 7.9290 0.4770 ;
      RECT 7.8790 0.1260 7.9290 0.4270 ;
      RECT 0.7190 0.5100 1.2570 0.5600 ;
      RECT 1.1750 1.1330 1.5610 1.1830 ;
      RECT 0.7190 0.9410 0.9530 0.9910 ;
      RECT 8.8510 1.1520 9.3890 1.2020 ;
      RECT 8.3190 0.2480 9.1610 0.2980 ;
      RECT 2.8630 0.7130 2.9890 0.7630 ;
      RECT 2.8630 0.7630 2.9130 1.0330 ;
      RECT 2.9390 0.5630 2.9890 0.7130 ;
      RECT 2.8470 0.5130 2.9890 0.5630 ;
      RECT 4.8230 0.3880 5.4970 0.4380 ;
      RECT 5.4470 0.4380 5.4970 0.5630 ;
      RECT 5.4470 0.2970 5.4970 0.3880 ;
      RECT 5.2950 0.9670 5.5130 1.0170 ;
      RECT 5.2950 0.3840 5.3450 0.3880 ;
    LAYER PO ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 5.8370 0.0660 5.8670 0.6910 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 3.1010 0.8400 3.1310 1.6060 ;
      RECT 5.8370 0.9390 5.8670 1.6060 ;
      RECT 5.5330 0.0660 5.5630 0.6370 ;
      RECT 3.1010 0.0660 3.1310 0.6370 ;
      RECT 9.3330 0.0660 9.3630 1.6060 ;
      RECT 3.7090 0.0660 3.7390 0.6910 ;
      RECT 5.0770 0.0660 5.1070 0.6910 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 9.6370 0.0660 9.6670 1.6060 ;
      RECT 4.7730 0.8920 4.8030 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 5.5330 0.8390 5.5630 1.6060 ;
      RECT 9.7890 0.0660 9.8190 1.6060 ;
      RECT 10.2450 0.0660 10.2750 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 9.9410 0.0660 9.9710 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 10.0930 0.0660 10.1230 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 4.7730 0.0660 4.8030 0.6910 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 3.7090 0.9390 3.7390 1.6060 ;
      RECT 7.3570 0.0670 7.3870 1.6050 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 5.0770 0.8390 5.1070 1.6060 ;
      RECT 9.4850 0.0660 9.5150 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
    LAYER NWELL ;
      RECT 7.7120 0.4910 9.7230 1.0830 ;
      RECT -0.1150 1.5430 10.6220 1.7730 ;
      RECT -0.1150 0.6790 7.2500 1.5430 ;
      RECT 10.3470 0.6790 10.6220 1.5430 ;
  END
END RSDFFNSRASRNX1_LVT

MACRO RDFFNSRASRX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.816 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 8.8160 1.7020 ;
        RECT 0.2790 1.1310 0.3290 1.6420 ;
        RECT 0.4480 1.2940 0.4980 1.6420 ;
        RECT 2.1430 1.2700 2.1930 1.6420 ;
        RECT 6.8550 1.4540 6.9050 1.6420 ;
        RECT 0.4480 1.2440 0.9530 1.2940 ;
        RECT 1.9340 1.2200 3.2330 1.2700 ;
        RECT 3.9270 1.4040 6.9050 1.4540 ;
        RECT 3.9270 1.2790 3.9770 1.4040 ;
        RECT 4.9910 0.9130 5.0410 1.4040 ;
        RECT 5.5990 1.0530 5.6490 1.4040 ;
        RECT 5.2950 0.9610 5.3450 1.4040 ;
        RECT 4.6870 0.9530 4.7370 1.4040 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 8.8160 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.2640 ;
        RECT 7.8790 0.0300 7.9290 0.4260 ;
        RECT 5.5990 0.0300 5.6490 0.2210 ;
        RECT 5.2950 0.0300 5.3450 0.3200 ;
        RECT 4.9910 0.0300 5.0410 0.4090 ;
        RECT 7.4230 0.0300 7.4730 0.1980 ;
        RECT 6.5110 0.0300 6.5610 0.4260 ;
        RECT 4.8630 0.0300 4.9130 0.2930 ;
        RECT 0.2790 0.2640 2.1530 0.3140 ;
        RECT 3.9110 0.2930 4.9130 0.3430 ;
        RECT 1.9510 0.3140 2.0010 0.5570 ;
        RECT 0.7350 0.3140 0.7850 0.5570 ;
        RECT 0.8870 0.3140 0.9370 0.5570 ;
        RECT 2.1030 0.3140 2.1530 0.5330 ;
        RECT 0.2790 0.3140 0.3290 0.4050 ;
        RECT 2.1030 0.2440 2.1530 0.2640 ;
        RECT 2.1030 0.1940 3.2330 0.2440 ;
        RECT 2.5590 0.2440 2.6090 0.3490 ;
    END
  END VSS

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.1550 0.8570 4.3110 0.9750 ;
        RECT 4.1550 0.9750 4.2050 1.0790 ;
        RECT 3.6230 1.0790 4.2050 1.1290 ;
        RECT 3.6230 1.1290 3.6730 1.3200 ;
        RECT 2.3310 1.3200 3.6730 1.3700 ;
        RECT 2.3310 1.3700 2.3810 1.4550 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6150 0.0880 4.6610 0.1380 ;
        RECT 1.6150 0.1380 1.7730 0.2100 ;
        RECT 4.6110 0.1380 4.6610 0.1700 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.4210 0.6630 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.0010 0.2490 8.1130 0.3590 ;
        RECT 8.0120 0.3590 8.0620 0.5270 ;
        RECT 7.7870 0.5270 8.0620 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4470 0.1490 5.4970 0.2710 ;
        RECT 5.4470 0.2710 6.1460 0.3210 ;
        RECT 6.0250 0.3210 6.1460 0.3600 ;
        RECT 6.0250 0.2500 6.1460 0.2710 ;
        RECT 6.0960 0.3600 6.1460 0.9330 ;
        RECT 5.4470 0.9330 6.1460 0.9830 ;
        RECT 5.4470 0.9830 5.4970 1.3270 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8330 0.7050 2.9890 0.7310 ;
        RECT 2.8330 0.7310 3.2930 0.7810 ;
        RECT 2.9390 0.5970 2.9890 0.7050 ;
        RECT 2.8330 0.7810 2.9890 0.8150 ;
        RECT 3.2430 0.7810 3.2930 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.4650 0.7250 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 6.4950 0.9420 8.1130 1.0020 ;
        RECT 8.0030 0.6900 8.1130 0.9420 ;
        RECT 7.8790 0.6270 7.9290 0.9420 ;
    END
  END VDDG

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8720 0.3990 5.9860 0.4020 ;
        RECT 5.1430 0.4020 5.9960 0.4520 ;
        RECT 5.1430 0.1490 5.1930 0.4020 ;
        RECT 5.8720 0.4520 5.9960 0.5120 ;
        RECT 5.9460 0.5120 5.9960 0.8330 ;
        RECT 5.1430 0.8330 5.9960 0.8830 ;
        RECT 5.1430 0.8830 5.1930 1.3190 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN
  OBS
    LAYER PO ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 2.9490 0.0660 2.9790 0.6910 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 1.8850 0.9390 1.9150 1.6060 ;
      RECT 5.8370 0.0670 5.8670 1.6050 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 3.2530 0.8390 3.2830 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 4.0130 0.0660 4.0430 0.6910 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 1.2770 0.8400 1.3070 1.6060 ;
      RECT 4.0130 0.9390 4.0430 1.6060 ;
      RECT 3.7090 0.0660 3.7390 0.6370 ;
      RECT 1.2770 0.0660 1.3070 0.6370 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
      RECT 1.8850 0.0660 1.9150 0.6910 ;
      RECT 3.2530 0.0660 3.2830 0.6910 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 2.9490 0.8920 2.9790 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 3.7090 0.8390 3.7390 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
    LAYER NWELL ;
      RECT 6.1920 0.4910 8.2030 1.0830 ;
      RECT -0.1150 1.5430 8.9380 1.7730 ;
      RECT -0.1150 0.6790 5.7300 1.5430 ;
      RECT 8.6630 0.6790 8.9380 1.5430 ;
    LAYER M1 ;
      RECT 1.0390 0.7130 1.1650 0.7630 ;
      RECT 1.0390 0.7630 1.0890 1.0330 ;
      RECT 1.1150 0.5630 1.1650 0.7130 ;
      RECT 1.0230 0.5130 1.1650 0.5630 ;
      RECT 2.9990 0.3940 3.6730 0.4440 ;
      RECT 3.6230 0.4440 3.6730 0.5630 ;
      RECT 3.6230 0.2970 3.6730 0.3940 ;
      RECT 3.4710 0.9670 3.6890 1.0170 ;
      RECT 3.4710 0.4440 3.5210 0.9670 ;
      RECT 3.4710 1.0170 3.5210 1.1200 ;
      RECT 3.4710 1.1700 3.5210 1.2700 ;
      RECT 2.9990 1.1200 3.5210 1.1700 ;
      RECT 2.3890 0.8580 2.5490 0.9080 ;
      RECT 2.3890 0.9080 2.4390 0.9680 ;
      RECT 1.8590 0.9680 2.4390 1.0180 ;
      RECT 1.3430 0.8540 2.2450 0.9040 ;
      RECT 1.3430 0.9040 1.3930 1.0590 ;
      RECT 1.3430 0.6130 1.3930 0.8540 ;
      RECT 1.3430 1.0590 1.7130 1.1090 ;
      RECT 1.3430 0.5630 1.5450 0.6130 ;
      RECT 1.3430 1.1090 1.3930 1.3370 ;
      RECT 1.4950 0.4070 1.5450 0.5630 ;
      RECT 1.3430 0.4130 1.3930 0.5630 ;
      RECT 4.7210 0.6320 5.2860 0.6820 ;
      RECT 4.1190 0.4500 4.1690 0.7290 ;
      RECT 4.1190 0.7290 4.4850 0.7790 ;
      RECT 4.4350 0.7790 4.4850 1.1790 ;
      RECT 4.7630 0.4500 4.8130 0.6320 ;
      RECT 3.7750 0.4000 4.8130 0.4500 ;
      RECT 3.7760 1.1790 4.4850 1.2290 ;
      RECT 3.7750 0.4500 3.8250 0.5630 ;
      RECT 3.7750 0.2970 3.8250 0.4000 ;
      RECT 3.7760 1.2290 3.8260 1.3530 ;
      RECT 2.6190 1.5200 3.3090 1.5700 ;
      RECT 3.0740 0.6130 3.3090 0.6630 ;
      RECT 3.3590 0.5440 3.4090 1.0200 ;
      RECT 2.8470 0.5170 3.4090 0.5440 ;
      RECT 2.8630 1.0200 3.4090 1.0700 ;
      RECT 2.8470 0.4940 3.4080 0.5170 ;
      RECT 2.5990 0.7880 2.6490 1.1200 ;
      RECT 1.5500 0.7380 2.6510 0.7880 ;
      RECT 2.4070 0.5050 2.4570 0.7380 ;
      RECT 2.8630 1.0700 2.9130 1.1200 ;
      RECT 2.0870 1.1200 2.9130 1.1700 ;
      RECT 3.6230 0.8670 3.7650 0.9170 ;
      RECT 3.6230 0.6630 3.6730 0.8670 ;
      RECT 3.6230 0.6130 4.0690 0.6630 ;
      RECT 2.7110 0.9200 3.1410 0.9700 ;
      RECT 3.0910 0.8310 3.1410 0.9200 ;
      RECT 2.7110 0.9700 2.7610 1.0340 ;
      RECT 2.7110 0.5050 2.7610 0.9200 ;
      RECT 2.4670 1.4200 3.7730 1.4700 ;
      RECT 1.4790 1.1900 1.8650 1.2400 ;
      RECT 4.0560 1.2870 4.4490 1.3370 ;
      RECT 1.4030 1.3890 1.9410 1.4390 ;
      RECT 3.3230 0.1880 3.9170 0.2380 ;
      RECT 3.3230 0.2380 3.3730 0.2940 ;
      RECT 2.6820 0.2940 3.3730 0.3440 ;
      RECT 2.2950 0.4550 2.3450 0.6130 ;
      RECT 1.8590 0.6130 2.3450 0.6630 ;
      RECT 2.6820 0.3440 2.7320 0.4050 ;
      RECT 2.2950 0.4050 2.7320 0.4550 ;
      RECT 0.7950 1.5240 2.0930 1.5740 ;
      RECT 1.1910 0.8130 1.2810 0.8630 ;
      RECT 1.1910 0.8630 1.2410 1.0830 ;
      RECT 1.2310 0.4620 1.2810 0.8130 ;
      RECT 0.4310 1.0830 1.2410 1.1330 ;
      RECT 1.1750 0.4120 1.2810 0.4620 ;
      RECT 1.1910 1.1330 1.2410 1.3540 ;
      RECT 0.4310 0.7980 0.4810 1.0830 ;
      RECT 0.4310 0.7480 0.5210 0.7980 ;
      RECT 0.4310 0.4350 0.5210 0.4850 ;
      RECT 0.4310 0.3720 0.4810 0.4350 ;
      RECT 0.4710 0.4850 0.5210 0.7480 ;
      RECT 5.3520 0.6130 5.8930 0.6630 ;
      RECT 4.5350 0.7830 4.5850 1.3010 ;
      RECT 4.5350 0.5500 4.5850 0.7330 ;
      RECT 4.3070 0.5000 4.5850 0.5500 ;
      RECT 4.3070 0.5500 4.3570 0.6790 ;
      RECT 4.8390 0.7830 4.8890 1.3010 ;
      RECT 5.3520 0.6630 5.4020 0.7330 ;
      RECT 4.5350 0.7330 5.4020 0.7830 ;
      RECT 5.8110 1.1990 7.1090 1.2490 ;
      RECT 3.9340 0.9670 4.0690 1.0170 ;
      RECT 3.9340 0.9160 3.9840 0.9670 ;
      RECT 3.8350 0.8660 3.9840 0.9160 ;
      RECT 0.5830 0.6130 1.0290 0.6630 ;
      RECT 0.5830 0.6630 0.6330 1.0040 ;
      RECT 0.5830 0.4130 0.6330 0.6130 ;
      RECT 6.7990 0.8200 7.3470 0.8700 ;
      RECT 7.1030 0.7090 7.6410 0.7590 ;
      RECT 7.7270 0.6770 7.7770 0.7680 ;
      RECT 7.6870 0.4270 7.7770 0.4620 ;
      RECT 7.7270 0.1260 7.7770 0.4270 ;
      RECT 7.6870 0.6270 7.7770 0.6770 ;
      RECT 7.6870 0.5120 7.7370 0.6270 ;
      RECT 7.4830 0.4770 7.7370 0.5120 ;
      RECT 7.4830 0.4620 7.7770 0.4770 ;
      RECT 7.1030 0.1320 7.3370 0.1820 ;
      RECT 6.3590 1.0620 6.8080 1.1120 ;
      RECT 6.3590 0.6770 6.4090 1.0620 ;
      RECT 6.3190 0.6270 6.4090 0.6770 ;
      RECT 6.3190 0.4770 6.3690 0.6270 ;
      RECT 6.3190 0.4270 6.4090 0.4770 ;
      RECT 6.3590 0.1260 6.4090 0.4270 ;
      RECT 6.4190 0.5270 7.0170 0.5770 ;
      RECT 6.6630 0.5770 6.7130 0.8840 ;
      RECT 6.6630 0.1260 6.7130 0.5270 ;
      RECT 6.9670 0.5770 7.0170 0.7700 ;
      RECT 6.9670 0.3480 7.0170 0.5270 ;
      RECT 7.3310 1.0620 7.8690 1.1120 ;
      RECT 6.7990 0.2480 7.6410 0.2980 ;
      RECT 3.3770 1.5200 6.8050 1.5700 ;
      RECT 1.0980 0.0940 1.4910 0.1440 ;
  END
END RDFFNSRASRX2_LVT

MACRO RDFFNSRASX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.512 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 8.5120 1.7020 ;
        RECT 0.2790 1.1310 0.3290 1.6420 ;
        RECT 0.4480 1.2940 0.4980 1.6420 ;
        RECT 2.1430 1.2700 2.1930 1.6420 ;
        RECT 6.5510 1.4540 6.6010 1.6420 ;
        RECT 0.4480 1.2440 0.9530 1.2940 ;
        RECT 1.9340 1.2200 3.2330 1.2700 ;
        RECT 3.9270 1.4040 6.6010 1.4540 ;
        RECT 3.9270 1.2790 3.9770 1.4040 ;
        RECT 5.1430 0.9590 5.1930 1.4040 ;
        RECT 4.6870 0.9530 4.7370 1.4040 ;
    END
  END VDD

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.9910 0.4010 5.6910 0.4510 ;
        RECT 4.9910 0.1570 5.0410 0.4010 ;
        RECT 5.5690 0.4510 5.6910 0.5380 ;
        RECT 5.6410 0.5380 5.6910 0.8590 ;
        RECT 4.9910 0.8590 5.6910 0.9090 ;
        RECT 4.9910 0.9090 5.0410 1.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2950 0.9690 5.8290 1.0190 ;
        RECT 5.7790 0.3510 5.8290 0.9690 ;
        RECT 5.2950 1.0190 5.5270 1.1290 ;
        RECT 5.2790 0.3010 5.8290 0.3510 ;
        RECT 5.2950 1.1290 5.3450 1.3270 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 8.5120 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.2720 ;
        RECT 5.1430 0.0300 5.1930 0.2410 ;
        RECT 7.1190 0.0300 7.1690 0.1980 ;
        RECT 7.5750 0.0300 7.6250 0.4260 ;
        RECT 6.2070 0.0300 6.2570 0.4260 ;
        RECT 4.8630 0.0300 4.9130 0.2880 ;
        RECT 0.2790 0.2720 2.1530 0.3220 ;
        RECT 3.9110 0.2880 4.9130 0.3380 ;
        RECT 1.9510 0.3220 2.0010 0.5570 ;
        RECT 0.7350 0.3220 0.7850 0.5570 ;
        RECT 0.8870 0.3220 0.9370 0.5570 ;
        RECT 2.1030 0.3220 2.1530 0.5330 ;
        RECT 0.2790 0.3220 0.3290 0.4050 ;
        RECT 2.1030 0.2380 2.1530 0.2720 ;
        RECT 2.1030 0.1880 3.2330 0.2380 ;
        RECT 2.5590 0.2380 2.6090 0.3490 ;
    END
  END VSS

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.1550 0.8570 4.3110 0.9750 ;
        RECT 4.1550 0.9750 4.2050 1.0790 ;
        RECT 3.6230 1.0790 4.2050 1.1290 ;
        RECT 3.6230 1.1290 3.6730 1.3200 ;
        RECT 2.3310 1.3200 3.6730 1.3700 ;
        RECT 2.3310 1.3700 2.3810 1.4550 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.4650 0.7250 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.4210 0.6630 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.6970 0.2490 7.8090 0.3590 ;
        RECT 7.7080 0.3590 7.7580 0.5270 ;
        RECT 7.4830 0.5270 7.7580 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8330 0.7050 2.9890 0.7310 ;
        RECT 2.8330 0.7310 3.2930 0.7810 ;
        RECT 2.9390 0.5970 2.9890 0.7050 ;
        RECT 2.8330 0.7810 2.9890 0.8150 ;
        RECT 3.2430 0.7810 3.2930 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 6.1910 0.9420 7.8090 1.0020 ;
        RECT 7.6990 0.6900 7.8090 0.9420 ;
        RECT 7.5750 0.6270 7.6250 0.9420 ;
    END
  END VDDG
  OBS
    LAYER PO ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 2.9490 0.0660 2.9790 0.6910 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 1.8850 0.9390 1.9150 1.6060 ;
      RECT 5.5330 0.0670 5.5630 1.6050 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 3.2530 0.8390 3.2830 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 4.0130 0.0660 4.0430 0.6910 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 1.2770 0.8400 1.3070 1.6060 ;
      RECT 4.0130 0.9390 4.0430 1.6060 ;
      RECT 3.7090 0.0660 3.7390 0.6370 ;
      RECT 1.2770 0.0660 1.3070 0.6370 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 1.8850 0.0660 1.9150 0.6910 ;
      RECT 3.2530 0.0660 3.2830 0.6910 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 2.9490 0.8920 2.9790 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 3.7090 0.8390 3.7390 1.6060 ;
    LAYER NWELL ;
      RECT 5.8880 0.4910 7.8990 1.0830 ;
      RECT -0.1150 1.5430 8.6330 1.7730 ;
      RECT -0.1150 0.6790 5.4260 1.5430 ;
      RECT 8.3590 0.6790 8.6330 1.5430 ;
    LAYER M1 ;
      RECT 1.1150 0.5630 1.1650 0.7130 ;
      RECT 1.0390 0.7130 1.1650 0.7630 ;
      RECT 1.0230 0.5130 1.1650 0.5630 ;
      RECT 1.0390 0.7630 1.0890 1.0330 ;
      RECT 2.9990 0.3880 3.6730 0.4380 ;
      RECT 3.6230 0.4380 3.6730 0.5630 ;
      RECT 3.6230 0.2970 3.6730 0.3880 ;
      RECT 3.4710 0.9670 3.6890 1.0170 ;
      RECT 3.4710 0.3840 3.5210 0.3880 ;
      RECT 3.4710 0.4380 3.5210 0.9670 ;
      RECT 3.4710 1.0170 3.5210 1.1200 ;
      RECT 3.4710 1.1700 3.5210 1.2700 ;
      RECT 2.9990 1.1200 3.5210 1.1700 ;
      RECT 2.3890 0.8580 2.5490 0.9080 ;
      RECT 2.3890 0.9080 2.4390 0.9680 ;
      RECT 1.8590 0.9680 2.4390 1.0180 ;
      RECT 1.3430 0.8540 2.2450 0.9040 ;
      RECT 1.3430 0.9040 1.3930 1.0590 ;
      RECT 1.3430 0.6130 1.3930 0.8540 ;
      RECT 1.3430 1.0590 1.7130 1.1090 ;
      RECT 1.3430 0.5630 1.5450 0.6130 ;
      RECT 1.3430 1.1090 1.3930 1.3370 ;
      RECT 1.4950 0.4070 1.5450 0.5630 ;
      RECT 1.3430 0.4130 1.3930 0.5630 ;
      RECT 4.7630 0.6420 5.1170 0.6920 ;
      RECT 5.0670 0.5970 5.1170 0.6420 ;
      RECT 4.1190 0.4500 4.1690 0.7290 ;
      RECT 4.1190 0.7290 4.4850 0.7790 ;
      RECT 4.4350 0.7790 4.4850 1.1790 ;
      RECT 4.7630 0.4500 4.8130 0.6420 ;
      RECT 3.7750 0.4000 4.8130 0.4500 ;
      RECT 3.7760 1.1790 4.4850 1.2290 ;
      RECT 3.7750 0.4500 3.8250 0.5630 ;
      RECT 3.7750 0.2970 3.8250 0.4000 ;
      RECT 3.7760 1.2290 3.8260 1.3530 ;
      RECT 4.0560 1.2790 4.4490 1.3290 ;
      RECT 1.4030 1.3890 1.9410 1.4390 ;
      RECT 3.3230 0.1880 3.9170 0.2380 ;
      RECT 3.3230 0.2380 3.3730 0.2880 ;
      RECT 2.6820 0.2880 3.3730 0.3380 ;
      RECT 2.2950 0.4550 2.3450 0.6130 ;
      RECT 1.8590 0.6130 2.3450 0.6630 ;
      RECT 2.6820 0.3380 2.7320 0.4050 ;
      RECT 2.2950 0.4050 2.7320 0.4550 ;
      RECT 1.1910 0.8130 1.2810 0.8630 ;
      RECT 1.1910 0.8630 1.2410 1.0830 ;
      RECT 1.2310 0.4620 1.2810 0.8130 ;
      RECT 0.4310 1.0830 1.2410 1.1330 ;
      RECT 1.1750 0.4120 1.2810 0.4620 ;
      RECT 1.1910 1.1330 1.2410 1.3540 ;
      RECT 0.4310 0.7980 0.4810 1.0830 ;
      RECT 0.4310 0.7480 0.5210 0.7980 ;
      RECT 0.4310 0.4350 0.5210 0.4850 ;
      RECT 0.4310 0.3720 0.4810 0.4350 ;
      RECT 0.4710 0.4850 0.5210 0.7480 ;
      RECT 5.1670 0.6130 5.5890 0.6630 ;
      RECT 4.5350 0.8090 4.5850 1.3010 ;
      RECT 4.5350 0.5500 4.5850 0.7590 ;
      RECT 4.3070 0.5000 4.5850 0.5500 ;
      RECT 4.3070 0.5500 4.3570 0.6790 ;
      RECT 4.8390 0.8090 4.8890 1.3010 ;
      RECT 5.1670 0.6630 5.2170 0.7590 ;
      RECT 4.5350 0.7590 5.2170 0.8090 ;
      RECT 5.5070 1.1990 6.8050 1.2490 ;
      RECT 3.6230 0.8670 3.7650 0.9170 ;
      RECT 3.6230 0.6630 3.6730 0.8670 ;
      RECT 3.6230 0.6130 4.0690 0.6630 ;
      RECT 3.9340 0.9670 4.0690 1.0170 ;
      RECT 3.9340 0.9160 3.9840 0.9670 ;
      RECT 3.8350 0.8660 3.9840 0.9160 ;
      RECT 2.8470 0.4880 3.4080 0.5070 ;
      RECT 2.8470 0.5070 3.4090 0.5380 ;
      RECT 3.3590 0.5380 3.4090 1.0200 ;
      RECT 2.8630 1.0200 3.4090 1.0700 ;
      RECT 2.5990 0.7880 2.6490 1.1200 ;
      RECT 1.5500 0.7380 2.6510 0.7880 ;
      RECT 2.4070 0.5050 2.4570 0.7380 ;
      RECT 2.8630 1.0700 2.9130 1.1200 ;
      RECT 2.0870 1.1200 2.9130 1.1700 ;
      RECT 0.5830 0.6130 1.0290 0.6630 ;
      RECT 0.5830 0.6630 0.6330 1.0040 ;
      RECT 0.5830 0.4130 0.6330 0.6130 ;
      RECT 4.6110 0.1380 4.6610 0.1700 ;
      RECT 1.7230 0.0880 4.6610 0.1380 ;
      RECT 1.7230 0.1380 1.7730 0.1700 ;
      RECT 6.4950 0.8200 7.0430 0.8700 ;
      RECT 6.7990 0.7090 7.3370 0.7590 ;
      RECT 7.4230 0.6770 7.4730 0.7680 ;
      RECT 7.3830 0.4270 7.4730 0.4620 ;
      RECT 7.4230 0.1260 7.4730 0.4270 ;
      RECT 7.3830 0.6270 7.4730 0.6770 ;
      RECT 7.3830 0.5120 7.4330 0.6270 ;
      RECT 7.1790 0.4770 7.4330 0.5120 ;
      RECT 7.1790 0.4620 7.4730 0.4770 ;
      RECT 6.7990 0.1320 7.0330 0.1820 ;
      RECT 6.0550 1.0620 6.5040 1.1120 ;
      RECT 6.0550 0.6770 6.1050 1.0620 ;
      RECT 6.0150 0.6270 6.1050 0.6770 ;
      RECT 6.0150 0.4770 6.0650 0.6270 ;
      RECT 6.0150 0.4270 6.1050 0.4770 ;
      RECT 6.0550 0.1260 6.1050 0.4270 ;
      RECT 1.0980 0.0940 1.4910 0.1440 ;
      RECT 6.1150 0.5270 6.7130 0.5770 ;
      RECT 6.3590 0.5770 6.4090 0.8910 ;
      RECT 6.3590 0.1260 6.4090 0.5270 ;
      RECT 6.6630 0.5770 6.7130 0.7700 ;
      RECT 6.6630 0.3480 6.7130 0.5270 ;
      RECT 0.7950 1.5240 2.0930 1.5740 ;
      RECT 7.0270 1.0620 7.5650 1.1120 ;
      RECT 6.4950 0.2480 7.3370 0.2980 ;
      RECT 3.3770 1.5200 6.5010 1.5700 ;
      RECT 2.6190 1.5200 3.3090 1.5700 ;
      RECT 3.0740 0.6130 3.3090 0.6630 ;
      RECT 2.7110 0.9200 3.1410 0.9700 ;
      RECT 3.0910 0.8310 3.1410 0.9200 ;
      RECT 2.7110 0.9700 2.7610 1.0340 ;
      RECT 2.7110 0.5050 2.7610 0.9200 ;
      RECT 2.4670 1.4200 3.7730 1.4700 ;
      RECT 1.4790 1.1900 1.8650 1.2400 ;
  END
END RDFFNSRASX1_LVT

MACRO RDFFNSRASX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.816 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 8.8160 1.7020 ;
        RECT 0.2790 1.1310 0.3290 1.6420 ;
        RECT 0.4480 1.2940 0.4980 1.6420 ;
        RECT 2.1430 1.2700 2.1930 1.6420 ;
        RECT 6.8550 1.4540 6.9050 1.6420 ;
        RECT 0.4480 1.2440 0.9530 1.2940 ;
        RECT 1.9340 1.2200 3.2330 1.2700 ;
        RECT 3.9270 1.4040 6.9050 1.4540 ;
        RECT 3.9270 1.2790 3.9770 1.4040 ;
        RECT 5.5990 1.0520 5.6490 1.4040 ;
        RECT 5.2950 0.9600 5.3450 1.4040 ;
        RECT 4.9910 0.9120 5.0410 1.4040 ;
        RECT 4.6870 0.9530 4.7370 1.4040 ;
    END
  END VDD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4470 0.1480 5.4970 0.2700 ;
        RECT 5.4470 0.2700 6.1450 0.3200 ;
        RECT 6.0240 0.3200 6.1450 0.3590 ;
        RECT 6.0240 0.2490 6.1450 0.2700 ;
        RECT 6.0950 0.3590 6.1450 0.9420 ;
        RECT 5.4470 0.9420 6.1450 0.9920 ;
        RECT 5.4470 0.9920 5.4970 1.3260 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 8.8160 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.2720 ;
        RECT 7.8790 0.0300 7.9290 0.4260 ;
        RECT 4.9910 0.0300 5.0410 0.4080 ;
        RECT 5.5990 0.0300 5.6490 0.2200 ;
        RECT 7.4230 0.0300 7.4730 0.1980 ;
        RECT 5.2950 0.0300 5.3450 0.3190 ;
        RECT 6.5110 0.0300 6.5610 0.4260 ;
        RECT 4.8630 0.0300 4.9130 0.2880 ;
        RECT 0.2790 0.2720 2.1530 0.3220 ;
        RECT 3.9110 0.2880 4.9130 0.3380 ;
        RECT 1.9510 0.3220 2.0010 0.5570 ;
        RECT 0.7350 0.3220 0.7850 0.5570 ;
        RECT 0.8870 0.3220 0.9370 0.5570 ;
        RECT 2.1030 0.3220 2.1530 0.5330 ;
        RECT 0.2790 0.3220 0.3290 0.4050 ;
        RECT 2.1030 0.2380 2.1530 0.2720 ;
        RECT 2.1030 0.1880 3.2330 0.2380 ;
        RECT 2.5590 0.2380 2.6090 0.3490 ;
    END
  END VSS

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.1550 0.8570 4.3110 0.9750 ;
        RECT 4.1550 0.9750 4.2050 1.0790 ;
        RECT 3.6230 1.0790 4.2050 1.1290 ;
        RECT 3.6230 1.1290 3.6730 1.3200 ;
        RECT 2.3310 1.3200 3.6730 1.3700 ;
        RECT 2.3310 1.3700 2.3810 1.4550 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.4650 0.7250 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.4210 0.6630 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.1430 0.1480 5.1930 0.4010 ;
        RECT 5.1430 0.4010 5.9950 0.4510 ;
        RECT 5.8730 0.4510 5.9950 0.5110 ;
        RECT 5.9450 0.5110 5.9950 0.8420 ;
        RECT 5.1430 0.8420 5.9950 0.8920 ;
        RECT 5.1430 0.8920 5.1930 1.3180 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.0010 0.2490 8.1130 0.3590 ;
        RECT 8.0120 0.3590 8.0620 0.5270 ;
        RECT 7.7870 0.5270 8.0620 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8330 0.7050 2.9890 0.7310 ;
        RECT 2.8330 0.7310 3.2930 0.7810 ;
        RECT 2.9390 0.5970 2.9890 0.7050 ;
        RECT 2.8330 0.7810 2.9890 0.8150 ;
        RECT 3.2430 0.7810 3.2930 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 6.4950 0.9420 8.1130 1.0020 ;
        RECT 8.0030 0.6900 8.1130 0.9420 ;
        RECT 7.8790 0.6270 7.9290 0.9420 ;
    END
  END VDDG
  OBS
    LAYER PO ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 2.9490 0.0660 2.9790 0.6910 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 1.8850 0.9390 1.9150 1.6060 ;
      RECT 5.8370 0.0670 5.8670 1.6050 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 3.2530 0.8390 3.2830 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 4.0130 0.0660 4.0430 0.6910 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 1.2770 0.8400 1.3070 1.6060 ;
      RECT 4.0130 0.9390 4.0430 1.6060 ;
      RECT 3.7090 0.0660 3.7390 0.6370 ;
      RECT 1.2770 0.0660 1.3070 0.6370 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 1.8850 0.0660 1.9150 0.6910 ;
      RECT 3.2530 0.0660 3.2830 0.6910 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 2.9490 0.8920 2.9790 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 3.7090 0.8390 3.7390 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
    LAYER NWELL ;
      RECT 6.1920 0.4910 8.2030 1.0830 ;
      RECT -0.1150 1.5430 8.9380 1.7730 ;
      RECT -0.1150 0.6790 5.7300 1.5430 ;
      RECT 8.6630 0.6790 8.9380 1.5430 ;
    LAYER M1 ;
      RECT 1.0390 0.7130 1.1650 0.7630 ;
      RECT 1.0390 0.7630 1.0890 1.0330 ;
      RECT 1.1150 0.5630 1.1650 0.7130 ;
      RECT 1.0230 0.5130 1.1650 0.5630 ;
      RECT 2.9990 0.3880 3.6730 0.4380 ;
      RECT 3.6230 0.4380 3.6730 0.5630 ;
      RECT 3.6230 0.2970 3.6730 0.3880 ;
      RECT 3.4710 0.9670 3.6890 1.0170 ;
      RECT 3.4710 0.4380 3.5210 0.9670 ;
      RECT 3.4710 1.0170 3.5210 1.1200 ;
      RECT 3.4710 1.1700 3.5210 1.2700 ;
      RECT 2.9990 1.1200 3.5210 1.1700 ;
      RECT 2.3890 0.8580 2.5490 0.9080 ;
      RECT 2.3890 0.9080 2.4390 0.9680 ;
      RECT 1.8590 0.9680 2.4390 1.0180 ;
      RECT 1.3430 0.8540 2.2450 0.9040 ;
      RECT 1.3430 0.9040 1.3930 1.0590 ;
      RECT 1.3430 0.6130 1.3930 0.8540 ;
      RECT 1.3430 1.0590 1.7130 1.1090 ;
      RECT 1.3430 0.5630 1.5450 0.6130 ;
      RECT 1.3430 1.1090 1.3930 1.3370 ;
      RECT 1.4950 0.4070 1.5450 0.5630 ;
      RECT 1.3430 0.4130 1.3930 0.5630 ;
      RECT 4.7630 0.6420 5.2850 0.6920 ;
      RECT 4.1190 0.4500 4.1690 0.7290 ;
      RECT 4.1190 0.7290 4.4850 0.7790 ;
      RECT 4.4350 0.7790 4.4850 1.1790 ;
      RECT 4.7630 0.4500 4.8130 0.6420 ;
      RECT 3.7750 0.4000 4.8130 0.4500 ;
      RECT 3.7760 1.1790 4.4850 1.2290 ;
      RECT 3.7750 0.4500 3.8250 0.5630 ;
      RECT 3.7750 0.2970 3.8250 0.4000 ;
      RECT 3.7760 1.2290 3.8260 1.3530 ;
      RECT 5.3490 0.6130 5.8930 0.6630 ;
      RECT 4.5350 0.7920 4.5850 1.3010 ;
      RECT 4.5350 0.5500 4.5850 0.7420 ;
      RECT 4.3070 0.5000 4.5850 0.5500 ;
      RECT 4.3070 0.5500 4.3570 0.6790 ;
      RECT 4.8390 0.7920 4.8890 1.3010 ;
      RECT 5.3490 0.6630 5.3990 0.7420 ;
      RECT 4.5350 0.7420 5.3990 0.7920 ;
      RECT 2.6190 1.5200 3.3090 1.5700 ;
      RECT 3.0740 0.6130 3.3090 0.6630 ;
      RECT 2.8470 0.4880 3.4090 0.5380 ;
      RECT 3.3590 0.5380 3.4090 1.0200 ;
      RECT 2.8630 1.0200 3.4090 1.0700 ;
      RECT 2.5990 0.7880 2.6490 1.1200 ;
      RECT 1.5500 0.7380 2.6510 0.7880 ;
      RECT 2.4070 0.5050 2.4570 0.7380 ;
      RECT 2.8630 1.0700 2.9130 1.1200 ;
      RECT 2.0870 1.1200 2.9130 1.1700 ;
      RECT 3.6230 0.8670 3.7650 0.9170 ;
      RECT 3.6230 0.6630 3.6730 0.8670 ;
      RECT 3.6230 0.6130 4.0690 0.6630 ;
      RECT 2.7110 0.9200 3.1410 0.9700 ;
      RECT 3.0910 0.8310 3.1410 0.9200 ;
      RECT 2.7110 0.9700 2.7610 1.0340 ;
      RECT 2.7110 0.5050 2.7610 0.9200 ;
      RECT 2.4670 1.4200 3.7730 1.4700 ;
      RECT 1.4790 1.1900 1.8650 1.2400 ;
      RECT 4.0560 1.2790 4.4490 1.3290 ;
      RECT 1.4030 1.3890 1.9410 1.4390 ;
      RECT 3.3230 0.1880 3.9170 0.2380 ;
      RECT 3.3230 0.2380 3.3730 0.2880 ;
      RECT 2.6820 0.2880 3.3730 0.3380 ;
      RECT 2.2950 0.4550 2.3450 0.6130 ;
      RECT 1.8590 0.6130 2.3450 0.6630 ;
      RECT 2.6820 0.3380 2.7320 0.4050 ;
      RECT 2.2950 0.4050 2.7320 0.4550 ;
      RECT 1.1910 0.8130 1.2810 0.8630 ;
      RECT 1.1910 0.8630 1.2410 1.0830 ;
      RECT 1.2310 0.4620 1.2810 0.8130 ;
      RECT 0.4310 1.0830 1.2410 1.1330 ;
      RECT 1.1750 0.4120 1.2810 0.4620 ;
      RECT 1.1910 1.1330 1.2410 1.3540 ;
      RECT 0.4310 0.7980 0.4810 1.0830 ;
      RECT 0.4310 0.7480 0.5210 0.7980 ;
      RECT 0.4310 0.4350 0.5210 0.4850 ;
      RECT 0.4310 0.3720 0.4810 0.4350 ;
      RECT 0.4710 0.4850 0.5210 0.7480 ;
      RECT 5.8110 1.1990 7.1090 1.2490 ;
      RECT 3.9340 0.9670 4.0690 1.0170 ;
      RECT 3.9340 0.9160 3.9840 0.9670 ;
      RECT 3.8350 0.8660 3.9840 0.9160 ;
      RECT 0.5830 0.6130 1.0290 0.6630 ;
      RECT 0.5830 0.6630 0.6330 1.0040 ;
      RECT 0.5830 0.4130 0.6330 0.6130 ;
      RECT 4.6110 0.1380 4.6610 0.1700 ;
      RECT 1.7230 0.0880 4.6610 0.1380 ;
      RECT 1.7230 0.1380 1.7730 0.1700 ;
      RECT 6.7990 0.8200 7.3470 0.8700 ;
      RECT 7.1030 0.7090 7.6410 0.7590 ;
      RECT 7.7270 0.6770 7.7770 0.7680 ;
      RECT 7.6870 0.4270 7.7770 0.4620 ;
      RECT 7.7270 0.1260 7.7770 0.4270 ;
      RECT 7.6870 0.6270 7.7770 0.6770 ;
      RECT 7.6870 0.5120 7.7370 0.6270 ;
      RECT 7.4830 0.4770 7.7370 0.5120 ;
      RECT 7.4830 0.4620 7.7770 0.4770 ;
      RECT 7.1030 0.1320 7.3370 0.1820 ;
      RECT 6.3590 1.0620 6.8080 1.1120 ;
      RECT 6.3590 0.6770 6.4090 1.0620 ;
      RECT 6.3190 0.6270 6.4090 0.6770 ;
      RECT 6.3190 0.4770 6.3690 0.6270 ;
      RECT 6.3190 0.4270 6.4090 0.4770 ;
      RECT 6.3590 0.1260 6.4090 0.4270 ;
      RECT 1.0980 0.0940 1.4910 0.1440 ;
      RECT 6.4190 0.5270 7.0170 0.5770 ;
      RECT 6.6630 0.5770 6.7130 0.8840 ;
      RECT 6.6630 0.1260 6.7130 0.5270 ;
      RECT 6.9670 0.5770 7.0170 0.7700 ;
      RECT 6.9670 0.3480 7.0170 0.5270 ;
      RECT 0.7950 1.5240 2.0930 1.5740 ;
      RECT 7.3310 1.0620 7.8690 1.1120 ;
      RECT 6.7990 0.2480 7.6410 0.2980 ;
      RECT 3.3770 1.5200 6.8050 1.5700 ;
  END
END RDFFNSRASX2_LVT

MACRO RDFFNSRX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.904 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 7.9040 1.7020 ;
        RECT 0.2790 1.1310 0.3290 1.6420 ;
        RECT 1.9910 1.2700 2.0410 1.6420 ;
        RECT 5.9430 1.4540 5.9930 1.6420 ;
        RECT 0.4480 1.2940 0.4980 1.6420 ;
        RECT 1.7830 1.2200 2.9290 1.2700 ;
        RECT 3.6230 1.4040 5.9930 1.4540 ;
        RECT 0.4480 1.2440 0.9530 1.2940 ;
        RECT 3.6230 1.2790 3.6730 1.4040 ;
        RECT 4.5350 0.9590 4.5850 1.4040 ;
        RECT 4.0790 0.9530 4.1290 1.4040 ;
    END
  END VDD

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.3830 0.4010 5.0830 0.4510 ;
        RECT 4.3830 0.1570 4.4330 0.4010 ;
        RECT 4.9610 0.4510 5.0830 0.5380 ;
        RECT 5.0330 0.5380 5.0830 0.8590 ;
        RECT 4.3830 0.8590 5.0830 0.9090 ;
        RECT 4.3830 0.9090 4.4330 1.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6870 0.9690 5.2210 1.0190 ;
        RECT 5.1710 0.3510 5.2210 0.9690 ;
        RECT 4.6870 1.0190 4.9190 1.1290 ;
        RECT 4.6710 0.3010 5.2210 0.3510 ;
        RECT 4.6870 1.1290 4.7370 1.3270 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.4650 0.7250 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 7.9040 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.2570 ;
        RECT 6.5110 0.0300 6.5610 0.1980 ;
        RECT 6.9670 0.0300 7.0170 0.4260 ;
        RECT 4.5350 0.0300 4.5850 0.2410 ;
        RECT 5.5990 0.0300 5.6490 0.4260 ;
        RECT 4.2550 0.0300 4.3050 0.2830 ;
        RECT 0.2790 0.2570 2.0010 0.3070 ;
        RECT 3.6070 0.2830 4.3050 0.3330 ;
        RECT 0.7350 0.3070 0.7850 0.5570 ;
        RECT 0.8870 0.3070 0.9370 0.5570 ;
        RECT 0.2790 0.3070 0.3290 0.4050 ;
        RECT 1.9510 0.2340 2.0010 0.2570 ;
        RECT 1.9510 0.1840 2.9290 0.2340 ;
        RECT 2.2550 0.2340 2.3050 0.3490 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.4210 0.6630 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.0850 0.2490 7.2010 0.3590 ;
        RECT 7.1000 0.3590 7.1500 0.5030 ;
        RECT 6.8750 0.5030 7.1500 0.5530 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5290 0.7050 2.6850 0.7310 ;
        RECT 2.5290 0.7310 2.9890 0.7810 ;
        RECT 2.6350 0.5970 2.6850 0.7050 ;
        RECT 2.5290 0.7810 2.6850 0.8150 ;
        RECT 2.9390 0.7810 2.9890 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 5.5830 0.9420 7.2010 1.0020 ;
        RECT 7.0910 0.6900 7.2010 0.9420 ;
        RECT 6.9670 0.6270 7.0170 0.9420 ;
    END
  END VDDG
  OBS
    LAYER PO ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 2.9490 0.8390 2.9790 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 1.7330 0.7300 1.7630 1.6060 ;
      RECT 3.7090 0.0660 3.7390 0.6910 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 1.2770 0.8400 1.3070 1.6060 ;
      RECT 3.7090 0.9390 3.7390 1.6060 ;
      RECT 3.4050 0.0660 3.4350 0.6370 ;
      RECT 1.2770 0.0660 1.3070 0.6370 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 2.9490 0.0660 2.9790 0.6910 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 2.6450 0.8920 2.6750 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 3.4050 0.8390 3.4350 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 1.7330 0.0680 1.7630 0.6180 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 2.6450 0.0660 2.6750 0.6910 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 4.9250 0.0670 4.9550 1.6050 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
    LAYER NWELL ;
      RECT 5.2800 0.4910 7.2910 1.0830 ;
      RECT -0.1150 1.5430 8.0260 1.7730 ;
      RECT -0.1150 0.6790 4.8180 1.5430 ;
      RECT 7.7510 0.6790 8.0260 1.5430 ;
    LAYER M1 ;
      RECT 4.1390 0.6320 4.5090 0.6820 ;
      RECT 4.4590 0.5970 4.5090 0.6320 ;
      RECT 3.8360 0.4500 3.8860 1.1790 ;
      RECT 3.4720 1.1790 3.9930 1.2290 ;
      RECT 4.2650 0.4500 4.3150 0.6320 ;
      RECT 3.4710 0.4000 4.3150 0.4500 ;
      RECT 3.4710 0.4500 3.5210 0.5630 ;
      RECT 3.4710 0.2970 3.5210 0.4000 ;
      RECT 3.4720 1.2290 3.5220 1.3530 ;
      RECT 4.8990 1.1990 6.1970 1.2490 ;
      RECT 0.4310 1.0830 1.2410 1.1330 ;
      RECT 1.1910 1.1330 1.2410 1.3540 ;
      RECT 1.1910 0.8630 1.2410 1.0830 ;
      RECT 1.1910 0.8130 1.2810 0.8630 ;
      RECT 1.2310 0.4620 1.2810 0.8130 ;
      RECT 1.1750 0.4120 1.2810 0.4620 ;
      RECT 0.4310 0.8690 0.4810 1.0830 ;
      RECT 0.4310 0.8190 0.5210 0.8690 ;
      RECT 0.4310 0.4250 0.5210 0.4750 ;
      RECT 0.4310 0.3620 0.4810 0.4250 ;
      RECT 0.4710 0.4750 0.5210 0.8190 ;
      RECT 3.3190 0.8670 3.4610 0.9170 ;
      RECT 3.3190 0.6630 3.3690 0.8670 ;
      RECT 3.3190 0.6130 3.7650 0.6630 ;
      RECT 3.0190 0.1780 3.6130 0.2280 ;
      RECT 3.0190 0.2280 3.0690 0.2840 ;
      RECT 2.3780 0.2840 3.0690 0.3340 ;
      RECT 1.7230 0.5240 1.7730 0.6130 ;
      RECT 1.9580 0.4550 2.0080 0.6130 ;
      RECT 1.7230 0.6130 2.0080 0.6630 ;
      RECT 2.3780 0.3340 2.4280 0.4050 ;
      RECT 1.9580 0.4050 2.4280 0.4550 ;
      RECT 3.6300 0.9670 3.7650 1.0170 ;
      RECT 3.6300 0.9160 3.6800 0.9670 ;
      RECT 3.5310 0.8660 3.6800 0.9160 ;
      RECT 2.5430 0.4840 3.1040 0.5070 ;
      RECT 2.5430 0.5070 3.1050 0.5340 ;
      RECT 3.0550 0.5340 3.1050 1.0200 ;
      RECT 2.5590 1.0200 3.1050 1.0700 ;
      RECT 2.2950 0.7880 2.3450 1.1200 ;
      RECT 1.5490 0.7380 2.3470 0.7880 ;
      RECT 2.1030 0.5050 2.1530 0.7380 ;
      RECT 2.5590 1.0700 2.6090 1.1200 ;
      RECT 1.9350 1.1200 2.6090 1.1700 ;
      RECT 4.5590 0.6130 4.9810 0.6630 ;
      RECT 4.0030 0.5670 4.0530 0.7590 ;
      RECT 4.2310 0.8090 4.2810 1.3010 ;
      RECT 4.0020 0.5170 4.1450 0.5670 ;
      RECT 4.5590 0.6630 4.6090 0.7590 ;
      RECT 4.0020 0.7590 4.6090 0.8090 ;
      RECT 0.5830 0.6130 1.0290 0.6630 ;
      RECT 0.5830 0.6630 0.6330 1.0040 ;
      RECT 0.5830 0.4130 0.6330 0.6130 ;
      RECT 1.0980 0.0940 1.4910 0.1440 ;
      RECT 5.8870 0.8200 6.4350 0.8700 ;
      RECT 1.3430 0.8540 2.0930 0.9040 ;
      RECT 1.3430 0.4840 1.3930 0.8540 ;
      RECT 1.3430 0.9040 1.3930 1.0990 ;
      RECT 1.3430 0.4340 1.5610 0.4840 ;
      RECT 1.3430 1.0990 1.5610 1.1490 ;
      RECT 1.3430 0.4080 1.3930 0.4340 ;
      RECT 1.3430 1.1490 1.3930 1.3370 ;
      RECT 6.1910 0.7090 6.7290 0.7590 ;
      RECT 1.4030 1.4240 1.7890 1.4740 ;
      RECT 6.7750 0.3920 6.8650 0.4420 ;
      RECT 6.7750 0.6270 6.8650 0.6770 ;
      RECT 6.8150 0.1260 6.8650 0.3920 ;
      RECT 6.8150 0.6770 6.8650 0.7680 ;
      RECT 6.5710 0.4620 6.8250 0.5120 ;
      RECT 6.7750 0.4420 6.8250 0.4620 ;
      RECT 6.7750 0.5120 6.8250 0.6270 ;
      RECT 6.1910 0.1320 6.4250 0.1820 ;
      RECT 5.4470 1.0770 5.8960 1.1270 ;
      RECT 5.4470 0.6770 5.4970 1.0770 ;
      RECT 5.4070 0.6270 5.4970 0.6770 ;
      RECT 5.4070 0.4770 5.4570 0.6270 ;
      RECT 5.4070 0.4270 5.4970 0.4770 ;
      RECT 5.4470 0.1260 5.4970 0.4270 ;
      RECT 0.7950 1.5240 1.9410 1.5740 ;
      RECT 5.5070 0.5270 6.1050 0.5770 ;
      RECT 5.7510 0.5770 5.8010 0.8770 ;
      RECT 5.7510 0.1260 5.8010 0.5270 ;
      RECT 6.0550 0.5770 6.1050 0.7700 ;
      RECT 6.0550 0.3480 6.1050 0.5270 ;
      RECT 3.8350 0.0960 4.0690 0.1460 ;
      RECT 6.4190 1.0860 6.9570 1.1360 ;
      RECT 5.8870 0.2480 6.7290 0.2980 ;
      RECT 3.0730 1.5200 5.8930 1.5700 ;
      RECT 2.3150 1.5200 3.0050 1.5700 ;
      RECT 2.7700 0.6130 3.0050 0.6630 ;
      RECT 2.4070 0.9200 2.8370 0.9700 ;
      RECT 2.7870 0.8310 2.8370 0.9200 ;
      RECT 2.4070 0.9700 2.4570 1.0340 ;
      RECT 2.4070 0.5050 2.4570 0.9200 ;
      RECT 2.1630 1.4200 3.4690 1.4700 ;
      RECT 1.0390 0.7130 1.1650 0.7630 ;
      RECT 1.0390 0.7630 1.0890 1.0330 ;
      RECT 1.1150 0.5630 1.1650 0.7130 ;
      RECT 1.0230 0.5130 1.1650 0.5630 ;
      RECT 2.6950 0.3840 3.3690 0.4340 ;
      RECT 3.3190 0.4340 3.3690 0.5630 ;
      RECT 3.3190 0.2970 3.3690 0.3840 ;
      RECT 3.1670 0.4340 3.2170 0.9670 ;
      RECT 3.1670 0.9670 3.3850 1.0170 ;
      RECT 3.1670 1.0170 3.2170 1.1200 ;
      RECT 3.1670 1.1700 3.2170 1.2700 ;
      RECT 2.6950 1.1200 3.2170 1.1700 ;
      RECT 1.7030 0.9680 2.2150 1.0180 ;
      RECT 2.1620 0.9080 2.2120 0.9680 ;
      RECT 2.1620 0.8580 2.2450 0.9080 ;
  END
END RDFFNSRX1_LVT

MACRO RDFFNSRX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.208 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 8.2080 1.7020 ;
        RECT 0.2790 1.1310 0.3290 1.6420 ;
        RECT 0.4480 1.2940 0.4980 1.6420 ;
        RECT 1.9910 1.2700 2.0410 1.6420 ;
        RECT 6.2470 1.4540 6.2970 1.6420 ;
        RECT 0.4480 1.2440 0.9530 1.2940 ;
        RECT 1.7830 1.2200 2.9290 1.2700 ;
        RECT 3.6230 1.4040 6.2970 1.4540 ;
        RECT 3.6230 1.2790 3.6730 1.4040 ;
        RECT 4.9910 1.0530 5.0410 1.4040 ;
        RECT 4.6870 0.9610 4.7370 1.4040 ;
        RECT 4.3830 0.9130 4.4330 1.4040 ;
        RECT 4.0790 0.9530 4.1290 1.4040 ;
    END
  END VDD

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.4650 0.7250 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 8.2080 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.2570 ;
        RECT 4.9910 0.0300 5.0410 0.2210 ;
        RECT 4.6870 0.0300 4.7370 0.3200 ;
        RECT 4.3830 0.0300 4.4330 0.4090 ;
        RECT 6.8150 0.0300 6.8650 0.1980 ;
        RECT 7.2710 0.0300 7.3210 0.4260 ;
        RECT 5.9030 0.0300 5.9530 0.4260 ;
        RECT 4.2550 0.0300 4.3050 0.2830 ;
        RECT 0.2790 0.2570 2.0010 0.3070 ;
        RECT 3.6070 0.2830 4.3050 0.3330 ;
        RECT 0.7350 0.3070 0.7850 0.5570 ;
        RECT 0.8870 0.3070 0.9370 0.5570 ;
        RECT 0.2790 0.3070 0.3290 0.4050 ;
        RECT 1.9510 0.2340 2.0010 0.2570 ;
        RECT 1.9510 0.1840 2.9290 0.2340 ;
        RECT 2.2550 0.2340 2.3050 0.3490 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.4210 0.6630 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2650 0.4010 5.3770 0.4020 ;
        RECT 4.5350 0.4020 5.3870 0.4520 ;
        RECT 4.5350 0.1490 4.5850 0.4020 ;
        RECT 5.2650 0.4520 5.3870 0.5120 ;
        RECT 5.3370 0.5120 5.3870 0.8330 ;
        RECT 4.5350 0.8330 5.3870 0.8830 ;
        RECT 4.5350 0.8830 4.5850 1.3190 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8390 0.1490 4.8890 0.2710 ;
        RECT 4.8390 0.2710 5.5370 0.3210 ;
        RECT 5.4160 0.3210 5.5370 0.3600 ;
        RECT 5.4160 0.2500 5.5370 0.2710 ;
        RECT 5.4870 0.3600 5.5370 0.9330 ;
        RECT 5.4160 0.2490 5.5290 0.2500 ;
        RECT 4.8390 0.9330 5.5370 0.9830 ;
        RECT 4.8390 0.9830 4.8890 1.3270 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.3930 0.2490 7.5050 0.3590 ;
        RECT 7.4040 0.3590 7.4540 0.5270 ;
        RECT 7.1790 0.5270 7.4540 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5290 0.7050 2.6850 0.7310 ;
        RECT 2.5290 0.7310 2.9890 0.7810 ;
        RECT 2.6350 0.5970 2.6850 0.7050 ;
        RECT 2.5290 0.7810 2.6850 0.8150 ;
        RECT 2.9390 0.7810 2.9890 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 5.8870 0.9420 7.5050 1.0020 ;
        RECT 7.3950 0.6900 7.5050 0.9420 ;
        RECT 7.2710 0.6270 7.3210 0.9420 ;
    END
  END VDDG
  OBS
    LAYER PO ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 2.9490 0.8390 2.9790 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 1.7330 0.7300 1.7630 1.6060 ;
      RECT 3.7090 0.0660 3.7390 0.6910 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 1.2770 0.8400 1.3070 1.6060 ;
      RECT 3.7090 0.9390 3.7390 1.6060 ;
      RECT 3.4050 0.0660 3.4350 0.6370 ;
      RECT 1.2770 0.0660 1.3070 0.6370 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 2.9490 0.0660 2.9790 0.6910 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 2.6450 0.8920 2.6750 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
      RECT 3.4050 0.8390 3.4350 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 1.7330 0.0680 1.7630 0.6180 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 2.6450 0.0660 2.6750 0.6910 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 5.2290 0.0670 5.2590 1.6050 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
    LAYER NWELL ;
      RECT 5.5840 0.4910 7.5950 1.0830 ;
      RECT -0.1150 1.5430 8.3290 1.7730 ;
      RECT -0.1150 0.6790 5.1220 1.5430 ;
      RECT 8.0550 0.6790 8.3290 1.5430 ;
    LAYER M1 ;
      RECT 4.1390 0.6320 4.6770 0.6820 ;
      RECT 3.4710 0.4500 3.5210 0.5630 ;
      RECT 3.4710 0.2970 3.5210 0.4000 ;
      RECT 3.4720 1.2290 3.5220 1.3530 ;
      RECT 3.8360 0.4500 3.8860 1.1790 ;
      RECT 3.4720 1.1790 3.9930 1.2290 ;
      RECT 3.4710 0.4000 4.3150 0.4500 ;
      RECT 4.2650 0.4500 4.3150 0.6320 ;
      RECT 1.0390 0.7130 1.1650 0.7630 ;
      RECT 1.0390 0.7630 1.0890 1.0330 ;
      RECT 1.1150 0.5630 1.1650 0.7130 ;
      RECT 1.0230 0.5130 1.1650 0.5630 ;
      RECT 2.6950 0.3840 3.3690 0.4340 ;
      RECT 3.3190 0.4340 3.3690 0.5630 ;
      RECT 3.3190 0.2970 3.3690 0.3840 ;
      RECT 3.1670 0.4340 3.2170 0.9670 ;
      RECT 3.1670 0.9670 3.3850 1.0170 ;
      RECT 3.1670 1.0170 3.2170 1.1200 ;
      RECT 3.1670 1.1700 3.2170 1.2700 ;
      RECT 2.6950 1.1200 3.2170 1.1700 ;
      RECT 1.7030 0.9680 2.2150 1.0180 ;
      RECT 2.1620 0.9080 2.2120 0.9680 ;
      RECT 2.1620 0.8580 2.2450 0.9080 ;
      RECT 3.0190 0.1780 3.6130 0.2280 ;
      RECT 3.0190 0.2280 3.0690 0.2840 ;
      RECT 2.3780 0.2840 3.0690 0.3340 ;
      RECT 1.7230 0.5240 1.7730 0.6130 ;
      RECT 1.9580 0.4550 2.0080 0.6130 ;
      RECT 1.7230 0.6130 2.0080 0.6630 ;
      RECT 2.3780 0.3340 2.4280 0.4050 ;
      RECT 1.9580 0.4050 2.4280 0.4550 ;
      RECT 2.4070 0.9200 2.8370 0.9700 ;
      RECT 2.7870 0.8310 2.8370 0.9200 ;
      RECT 2.4070 0.9700 2.4570 1.0340 ;
      RECT 2.4070 0.5050 2.4570 0.9200 ;
      RECT 2.1630 1.4200 3.4690 1.4700 ;
      RECT 1.1910 0.8130 1.2810 0.8630 ;
      RECT 1.1910 0.8630 1.2410 1.0830 ;
      RECT 1.2310 0.4620 1.2810 0.8130 ;
      RECT 0.4310 1.0830 1.2410 1.1330 ;
      RECT 1.1750 0.4120 1.2810 0.4620 ;
      RECT 1.1910 1.1330 1.2410 1.3540 ;
      RECT 0.4310 0.8690 0.4810 1.0830 ;
      RECT 0.4310 0.8190 0.5210 0.8690 ;
      RECT 0.4310 0.4250 0.5210 0.4750 ;
      RECT 0.4310 0.3620 0.4810 0.4250 ;
      RECT 0.4710 0.4750 0.5210 0.8190 ;
      RECT 4.7370 0.6130 5.2850 0.6630 ;
      RECT 4.0030 0.7820 4.0530 0.8090 ;
      RECT 4.0030 0.5670 4.0530 0.7320 ;
      RECT 4.2310 0.7820 4.2810 1.3010 ;
      RECT 4.0020 0.5170 4.1450 0.5670 ;
      RECT 4.7370 0.6630 4.7870 0.7320 ;
      RECT 4.0020 0.7320 4.7870 0.7820 ;
      RECT 5.2030 1.1990 6.5010 1.2490 ;
      RECT 3.3190 0.8670 3.4610 0.9170 ;
      RECT 3.3190 0.6630 3.3690 0.8670 ;
      RECT 3.3190 0.6130 3.7650 0.6630 ;
      RECT 3.6300 0.9670 3.7650 1.0170 ;
      RECT 3.6300 0.9160 3.6800 0.9670 ;
      RECT 3.5310 0.8660 3.6800 0.9160 ;
      RECT 2.5430 0.4840 3.1040 0.5070 ;
      RECT 2.5430 0.5070 3.1050 0.5340 ;
      RECT 3.0550 0.5340 3.1050 1.0200 ;
      RECT 2.5590 1.0200 3.1050 1.0700 ;
      RECT 2.2950 0.7880 2.3450 1.1200 ;
      RECT 1.5490 0.7380 2.3470 0.7880 ;
      RECT 2.1030 0.5050 2.1530 0.7380 ;
      RECT 2.5590 1.0700 2.6090 1.1200 ;
      RECT 1.9350 1.1200 2.6090 1.1700 ;
      RECT 0.5830 0.6130 1.0290 0.6630 ;
      RECT 0.5830 0.6630 0.6330 1.0040 ;
      RECT 0.5830 0.4130 0.6330 0.6130 ;
      RECT 1.0980 0.0940 1.4910 0.1440 ;
      RECT 6.1910 0.8200 6.7390 0.8700 ;
      RECT 1.3430 0.8540 2.0930 0.9040 ;
      RECT 1.3430 0.4840 1.3930 0.8540 ;
      RECT 1.3430 0.9040 1.3930 1.0990 ;
      RECT 1.3430 0.4340 1.5610 0.4840 ;
      RECT 1.3430 1.0990 1.5610 1.1490 ;
      RECT 1.3430 0.4080 1.3930 0.4340 ;
      RECT 1.3430 1.1490 1.3930 1.3370 ;
      RECT 6.4950 0.7090 7.0330 0.7590 ;
      RECT 1.4030 1.4240 1.7890 1.4740 ;
      RECT 7.1190 0.6770 7.1690 0.7680 ;
      RECT 7.0790 0.4270 7.1690 0.4620 ;
      RECT 7.1190 0.1260 7.1690 0.4270 ;
      RECT 7.0790 0.6270 7.1690 0.6770 ;
      RECT 7.0790 0.5120 7.1290 0.6270 ;
      RECT 6.8750 0.4770 7.1290 0.5120 ;
      RECT 6.8750 0.4620 7.1690 0.4770 ;
      RECT 6.4950 0.1320 6.7290 0.1820 ;
      RECT 5.7510 1.0620 6.2000 1.1120 ;
      RECT 5.7510 0.6770 5.8010 1.0620 ;
      RECT 5.7110 0.6270 5.8010 0.6770 ;
      RECT 5.7110 0.4770 5.7610 0.6270 ;
      RECT 5.7110 0.4270 5.8010 0.4770 ;
      RECT 5.7510 0.1260 5.8010 0.4270 ;
      RECT 0.7950 1.5240 1.9410 1.5740 ;
      RECT 5.8110 0.5270 6.4090 0.5770 ;
      RECT 6.0550 0.5770 6.1050 0.8840 ;
      RECT 6.0550 0.1260 6.1050 0.5270 ;
      RECT 6.3590 0.5770 6.4090 0.7700 ;
      RECT 6.3590 0.3480 6.4090 0.5270 ;
      RECT 3.8350 0.0880 4.0690 0.1380 ;
      RECT 6.7230 1.0620 7.2610 1.1120 ;
      RECT 6.1910 0.2480 7.0330 0.2980 ;
      RECT 3.0730 1.5200 6.1970 1.5700 ;
      RECT 2.3150 1.5200 3.0050 1.5700 ;
      RECT 2.7700 0.6130 3.0050 0.6630 ;
  END
END RDFFNSRX2_LVT

MACRO RDFFNX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.36 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 6.1910 0.9420 7.6580 1.0020 ;
        RECT 7.5480 0.6900 7.6580 0.9420 ;
    END
  END VDDG

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 8.3600 0.0300 ;
        RECT 0.3840 0.0300 0.4340 0.3070 ;
        RECT 7.2710 0.0300 7.3210 0.3120 ;
        RECT 5.1430 0.0300 5.1930 0.2410 ;
        RECT 6.9670 0.0300 7.0170 0.2020 ;
        RECT 6.2070 0.0300 6.2570 0.2060 ;
        RECT 4.8790 0.0300 4.9290 0.2830 ;
        RECT 0.3840 0.3070 2.1530 0.3570 ;
        RECT 2.9990 0.2830 4.9300 0.3330 ;
        RECT 0.4310 0.3570 0.4810 0.5570 ;
        RECT 1.4950 0.3570 1.5450 0.5580 ;
        RECT 1.6470 0.3570 1.6970 0.5580 ;
        RECT 2.1030 0.3570 2.1530 0.5770 ;
        RECT 4.8390 0.3330 4.8890 0.4430 ;
    END
  END VSS

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 1.4650 0.4220 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2950 0.9690 5.8290 1.0190 ;
        RECT 5.7790 0.3510 5.8290 0.9690 ;
        RECT 5.2950 1.0190 5.5270 1.1290 ;
        RECT 5.2790 0.3010 5.8290 0.3510 ;
        RECT 5.2950 1.1290 5.3450 1.3270 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.9910 0.1570 5.0410 0.4010 ;
        RECT 4.9910 0.4010 5.6910 0.4510 ;
        RECT 5.5690 0.4510 5.6910 0.5380 ;
        RECT 5.6410 0.5380 5.6910 0.8590 ;
        RECT 4.9910 0.8590 5.6910 0.9090 ;
        RECT 4.9910 0.9090 5.0410 1.2320 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 8.3600 1.7020 ;
        RECT 0.1380 1.3400 0.1880 1.6420 ;
        RECT 3.2070 1.3400 3.2570 1.6420 ;
        RECT 0.1380 1.2900 5.1940 1.3400 ;
        RECT 3.0150 0.9730 3.0650 1.2900 ;
        RECT 5.1430 0.9590 5.1930 1.2900 ;
    END
  END VDD

  PIN RETN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.5130 1.4080 6.8980 1.4580 ;
        RECT 6.7850 1.3130 6.8980 1.4080 ;
    END
    ANTENNAGATEAREA 0.084 ;
  END RETN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0950 0.9670 1.1810 1.0170 ;
        RECT 0.0950 1.0170 0.2080 1.1190 ;
    END
    ANTENNAGATEAREA 0.018 ;
  END D
  OBS
    LAYER PO ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 3.5570 0.9590 3.5870 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 5.5330 0.0670 5.5630 1.6050 ;
      RECT 1.7330 0.9390 1.7630 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 1.7330 0.0660 1.7630 0.6370 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 0.9730 0.0660 1.0030 0.6910 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 2.1890 0.9390 2.2190 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 3.5570 0.0660 3.5870 0.6910 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 4.0130 0.0660 4.0430 0.7910 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 2.6450 0.0660 2.6750 0.6910 ;
      RECT 2.1890 0.0660 2.2190 0.6370 ;
      RECT 0.9730 0.8390 1.0030 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 4.0130 0.9390 4.0430 1.6060 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 2.6450 0.8390 2.6750 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 3.7090 0.0660 3.7390 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
    LAYER NWELL ;
      RECT -0.1160 1.5430 8.4700 1.7730 ;
      RECT -0.1160 0.6790 5.4270 1.5430 ;
      RECT 8.1950 0.6790 8.4700 1.5430 ;
      RECT 5.8890 0.4910 7.7350 1.0830 ;
    LAYER M1 ;
      RECT 7.1190 0.5890 7.3120 0.6390 ;
      RECT 7.2620 0.5120 7.3120 0.5890 ;
      RECT 7.2620 0.4620 7.4130 0.5120 ;
      RECT 7.2620 0.4120 7.3120 0.4620 ;
      RECT 7.1190 0.3620 7.3120 0.4120 ;
      RECT 7.1190 0.6390 7.1690 0.7820 ;
      RECT 7.1190 0.1260 7.1690 0.3620 ;
      RECT 2.8230 0.7670 2.9530 0.8170 ;
      RECT 2.9030 0.5630 2.9530 0.7670 ;
      RECT 2.8630 0.5130 2.9530 0.5630 ;
      RECT 2.7110 1.1900 2.9130 1.2400 ;
      RECT 2.7110 0.9740 2.7610 1.1900 ;
      RECT 2.8630 1.0240 2.9130 1.1900 ;
      RECT 2.8230 0.9740 2.9130 1.0240 ;
      RECT 2.8230 0.8170 2.8730 0.9740 ;
      RECT 2.8630 0.3270 2.9130 0.5130 ;
      RECT 2.7110 0.2770 2.9130 0.3270 ;
      RECT 2.7110 0.3270 2.7610 0.5560 ;
      RECT 0.7950 1.5240 2.8530 1.5740 ;
      RECT 0.4910 0.0940 2.5490 0.1440 ;
      RECT 3.1270 0.7670 3.3690 0.8170 ;
      RECT 3.3190 0.8170 3.3690 1.2400 ;
      RECT 3.1270 0.4530 3.1770 0.7670 ;
      RECT 3.0030 0.4030 3.3700 0.4530 ;
      RECT 3.3190 0.4530 3.3690 0.5770 ;
      RECT 3.0030 0.4530 3.0530 0.8670 ;
      RECT 2.9230 0.8670 3.0530 0.9170 ;
      RECT 3.4310 0.5130 4.2970 0.5630 ;
      RECT 3.4310 0.5630 3.4810 0.6270 ;
      RECT 3.2270 0.6270 3.4810 0.6770 ;
      RECT 3.4310 0.6770 3.4810 1.0670 ;
      RECT 3.4310 1.0670 4.2970 1.1170 ;
      RECT 3.5310 0.6130 4.4330 0.6630 ;
      RECT 4.3830 0.3830 4.4330 0.6130 ;
      RECT 3.7350 0.6630 3.7850 0.9670 ;
      RECT 3.7350 0.9670 4.4330 1.0170 ;
      RECT 4.3830 1.0170 4.4330 1.2400 ;
      RECT 6.8150 0.4620 7.1090 0.5120 ;
      RECT 6.8150 0.1820 6.8650 0.4620 ;
      RECT 6.8150 0.5120 6.8650 0.6350 ;
      RECT 6.4950 0.1320 6.8650 0.1820 ;
      RECT 6.4950 0.6350 6.8650 0.6850 ;
      RECT 6.3590 0.4940 6.7130 0.5440 ;
      RECT 6.6630 0.3480 6.7130 0.4940 ;
      RECT 6.3590 0.5440 6.4090 0.7820 ;
      RECT 4.1390 0.7590 5.5890 0.8090 ;
      RECT 5.0670 0.6420 5.1170 0.7590 ;
      RECT 4.6870 0.8090 4.7370 1.2400 ;
      RECT 4.4950 0.5630 4.5450 0.7590 ;
      RECT 4.4950 0.5130 4.7370 0.5630 ;
      RECT 4.6870 0.3830 4.7370 0.5130 ;
      RECT 3.6830 1.5280 7.7190 1.5780 ;
      RECT 3.8350 0.7130 4.0690 0.7630 ;
      RECT 1.4790 0.9670 2.0930 1.0170 ;
      RECT 1.3430 0.4070 1.3930 0.6190 ;
      RECT 1.6470 0.6690 1.6970 0.9670 ;
      RECT 1.3430 0.6190 1.6970 0.6690 ;
      RECT 7.4230 0.5620 7.7170 0.6120 ;
      RECT 7.5580 0.4120 7.6080 0.5620 ;
      RECT 7.4230 0.3620 7.6080 0.4120 ;
      RECT 7.4230 0.6120 7.4730 0.8320 ;
      RECT 6.2590 0.8320 7.4730 0.8820 ;
      RECT 7.4230 0.1260 7.4730 0.3620 ;
      RECT 6.2590 0.4200 6.3090 0.8320 ;
      RECT 6.2590 0.3700 6.4270 0.4200 ;
      RECT 2.4670 0.8670 2.7210 0.9170 ;
      RECT 0.2790 0.6130 0.7250 0.6630 ;
      RECT 0.2790 0.8670 1.0290 0.9170 ;
      RECT 0.2790 0.4130 0.3290 0.6130 ;
      RECT 0.2790 0.6630 0.3290 0.8670 ;
      RECT 0.7190 0.5130 0.8610 0.5630 ;
      RECT 0.8110 0.5630 0.8610 0.6130 ;
      RECT 0.8110 0.6130 1.0290 0.6630 ;
      RECT 0.8110 0.6630 0.8610 0.7540 ;
      RECT 0.7180 0.7540 0.8610 0.8040 ;
      RECT 1.9110 0.8670 2.1930 0.9170 ;
      RECT 2.1430 0.9170 2.1930 1.1270 ;
      RECT 1.1910 1.1270 2.1930 1.1770 ;
      RECT 1.1910 1.1770 1.2410 1.2400 ;
      RECT 1.2410 0.9170 1.2910 1.0660 ;
      RECT 1.1910 0.4130 1.2410 0.8670 ;
      RECT 1.9110 0.6070 1.9610 0.8670 ;
      RECT 1.9110 0.5570 2.0010 0.6070 ;
      RECT 1.9510 0.4130 2.0010 0.5570 ;
      RECT 1.1910 1.0670 1.2910 1.1270 ;
      RECT 1.2310 1.0660 1.2910 1.0670 ;
      RECT 1.1910 0.8670 1.4850 0.9170 ;
      RECT 2.0110 0.6670 2.3970 0.7170 ;
      RECT 5.5070 1.2000 6.6530 1.2500 ;
      RECT 2.6190 0.6130 2.8530 0.6630 ;
      RECT 4.9670 0.5010 5.2690 0.5510 ;
      RECT 5.2190 0.5510 5.2690 0.6790 ;
      RECT 4.9670 0.5510 5.0170 0.6130 ;
      RECT 4.5950 0.6130 5.0170 0.6630 ;
      RECT 6.0550 1.0620 6.5010 1.1120 ;
      RECT 6.0550 0.1260 6.1050 1.0620 ;
      RECT 2.5990 0.0920 4.6780 0.1420 ;
      RECT 2.5990 0.1420 2.6490 0.1940 ;
      RECT 2.5590 0.1940 2.6490 0.2440 ;
      RECT 2.5590 0.2440 2.6090 0.5130 ;
      RECT 2.4070 0.5130 2.6090 0.5630 ;
      RECT 2.4070 0.2770 2.4570 0.5130 ;
      RECT 2.4470 0.5630 2.4970 0.7670 ;
      RECT 2.3670 0.7670 2.4970 0.8170 ;
      RECT 2.3670 0.8170 2.4170 0.9670 ;
      RECT 2.3670 0.9670 2.4570 1.0170 ;
      RECT 2.4070 1.0170 2.4570 1.1900 ;
      RECT 2.4070 1.1900 2.6090 1.2400 ;
      RECT 2.5590 0.9740 2.6090 1.1900 ;
  END
END RDFFNX1_LVT

MACRO RDFFNX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.664 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 6.4950 0.9420 7.9620 1.0020 ;
        RECT 7.8520 0.6900 7.9620 0.9420 ;
    END
  END VDDG

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.0250 0.3210 6.1450 0.3600 ;
        RECT 5.4470 0.2710 6.1450 0.3210 ;
        RECT 6.0950 0.3600 6.1450 0.9330 ;
        RECT 6.0250 0.2500 6.1450 0.2710 ;
        RECT 5.4470 0.1490 5.4970 0.2710 ;
        RECT 5.4470 0.9330 6.1450 0.9830 ;
        RECT 6.0250 0.2490 6.1370 0.2500 ;
        RECT 5.4470 0.9830 5.4970 1.2240 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8730 0.4000 5.9850 0.4020 ;
        RECT 5.1430 0.4020 5.9950 0.4520 ;
        RECT 5.1430 0.1490 5.1930 0.4020 ;
        RECT 5.8730 0.4520 5.9950 0.5120 ;
        RECT 5.9450 0.5120 5.9950 0.8330 ;
        RECT 5.1430 0.8330 5.9950 0.8830 ;
        RECT 5.1430 0.8830 5.1930 1.2240 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 8.6640 0.0300 ;
        RECT 0.3840 0.0300 0.4340 0.3070 ;
        RECT 7.5750 0.0300 7.6250 0.3120 ;
        RECT 6.5110 0.0300 6.5610 0.2060 ;
        RECT 5.2950 0.0300 5.3450 0.3200 ;
        RECT 7.2710 0.0300 7.3210 0.2020 ;
        RECT 5.5990 0.0300 5.6490 0.2210 ;
        RECT 4.9910 0.0300 5.0410 0.4090 ;
        RECT 4.8790 0.0300 4.9290 0.2830 ;
        RECT 0.3840 0.3070 2.1530 0.3570 ;
        RECT 2.9990 0.2830 4.9300 0.3330 ;
        RECT 0.4310 0.3570 0.4810 0.5570 ;
        RECT 2.1030 0.3570 2.1530 0.5770 ;
        RECT 1.4950 0.3570 1.5450 0.5580 ;
        RECT 1.6470 0.3570 1.6970 0.5580 ;
        RECT 4.8390 0.3330 4.8890 0.4430 ;
    END
  END VSS

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2480 1.4650 0.4220 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 8.6640 1.7020 ;
        RECT 0.1380 1.3400 0.1880 1.6420 ;
        RECT 3.2070 1.3400 3.2570 1.6420 ;
        RECT 0.1380 1.2900 5.6490 1.3400 ;
        RECT 5.5990 1.0530 5.6490 1.2900 ;
        RECT 4.9910 0.9130 5.0410 1.2900 ;
        RECT 5.2950 0.9610 5.3450 1.2900 ;
        RECT 3.0150 0.9730 3.0650 1.2900 ;
    END
  END VDD

  PIN RETN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.5130 1.4080 7.2020 1.4580 ;
        RECT 7.0890 1.3130 7.2020 1.4080 ;
    END
    ANTENNAGATEAREA 0.084 ;
  END RETN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0940 0.9670 1.1810 1.0170 ;
        RECT 0.0940 1.0170 0.2080 1.1190 ;
    END
    ANTENNAGATEAREA 0.018 ;
  END D
  OBS
    LAYER PO ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 3.5570 0.9590 3.5870 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 5.8370 0.0670 5.8670 1.6050 ;
      RECT 1.7330 0.9390 1.7630 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 1.7330 0.0660 1.7630 0.6370 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 0.9730 0.0660 1.0030 0.6910 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 2.1890 0.9390 2.2190 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 3.5570 0.0660 3.5870 0.6910 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 4.0130 0.0660 4.0430 0.7910 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 2.6450 0.0660 2.6750 0.6910 ;
      RECT 2.1890 0.0660 2.2190 0.6370 ;
      RECT 0.9730 0.8390 1.0030 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 4.0130 0.9390 4.0430 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 2.6450 0.8390 2.6750 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 3.7090 0.0660 3.7390 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
    LAYER NWELL ;
      RECT -0.1160 1.5430 8.7740 1.7730 ;
      RECT -0.1160 0.6790 5.7310 1.5430 ;
      RECT 8.4990 0.6790 8.7740 1.5430 ;
      RECT 6.1930 0.4910 8.0390 1.0830 ;
    LAYER M1 ;
      RECT 2.5990 0.0920 4.6780 0.1420 ;
      RECT 2.4070 1.0170 2.4570 1.1900 ;
      RECT 2.3670 0.9670 2.4570 1.0170 ;
      RECT 2.4070 1.1900 2.6090 1.2400 ;
      RECT 2.3670 0.8170 2.4170 0.9670 ;
      RECT 2.5590 0.9740 2.6090 1.1900 ;
      RECT 2.3670 0.7670 2.4970 0.8170 ;
      RECT 2.4470 0.5630 2.4970 0.7670 ;
      RECT 2.4070 0.5130 2.6090 0.5630 ;
      RECT 2.4070 0.2770 2.4570 0.5130 ;
      RECT 2.5590 0.2440 2.6090 0.5130 ;
      RECT 2.5590 0.1940 2.6490 0.2440 ;
      RECT 2.5990 0.1420 2.6490 0.1940 ;
      RECT 4.9180 0.5200 5.4030 0.5700 ;
      RECT 5.3530 0.5700 5.4030 0.6040 ;
      RECT 4.9180 0.5700 4.9680 0.6130 ;
      RECT 5.3530 0.6040 5.5890 0.6540 ;
      RECT 4.5950 0.6130 4.9680 0.6630 ;
      RECT 7.4230 0.5890 7.6160 0.6390 ;
      RECT 7.5660 0.5120 7.6160 0.5890 ;
      RECT 7.5660 0.4620 7.7170 0.5120 ;
      RECT 7.5660 0.4120 7.6160 0.4620 ;
      RECT 7.4230 0.3620 7.6160 0.4120 ;
      RECT 7.4230 0.6390 7.4730 0.7820 ;
      RECT 7.4230 0.1260 7.4730 0.3620 ;
      RECT 2.6190 0.6130 2.8530 0.6630 ;
      RECT 1.9110 0.8670 2.1930 0.9170 ;
      RECT 2.1430 0.9170 2.1930 1.1270 ;
      RECT 1.1910 1.1270 2.1930 1.1770 ;
      RECT 1.1910 1.1770 1.2410 1.2400 ;
      RECT 1.2410 0.9170 1.2910 1.0660 ;
      RECT 1.1910 0.4130 1.2410 0.8670 ;
      RECT 1.9110 0.6070 1.9610 0.8670 ;
      RECT 1.9110 0.5570 2.0010 0.6070 ;
      RECT 1.9510 0.4130 2.0010 0.5570 ;
      RECT 1.1910 1.0670 1.2910 1.1270 ;
      RECT 1.2310 1.0660 1.2910 1.0670 ;
      RECT 1.1910 0.8670 1.4850 0.9170 ;
      RECT 2.8230 0.7670 2.9530 0.8170 ;
      RECT 2.9030 0.5630 2.9530 0.7670 ;
      RECT 2.8630 0.5130 2.9530 0.5630 ;
      RECT 2.7110 1.1900 2.9130 1.2400 ;
      RECT 2.7110 0.9740 2.7610 1.1900 ;
      RECT 2.8630 1.0240 2.9130 1.1900 ;
      RECT 2.8230 0.9740 2.9130 1.0240 ;
      RECT 2.8230 0.8170 2.8730 0.9740 ;
      RECT 2.8630 0.3270 2.9130 0.5130 ;
      RECT 2.7110 0.2770 2.9130 0.3270 ;
      RECT 2.7110 0.3270 2.7610 0.5560 ;
      RECT 0.7950 1.5240 2.8530 1.5740 ;
      RECT 0.4910 0.0940 2.5490 0.1440 ;
      RECT 3.1270 0.7670 3.3690 0.8170 ;
      RECT 3.3190 0.8170 3.3690 1.2400 ;
      RECT 3.1270 0.4530 3.1770 0.7670 ;
      RECT 3.0030 0.4030 3.3700 0.4530 ;
      RECT 3.3190 0.4530 3.3690 0.5770 ;
      RECT 3.0030 0.4530 3.0530 0.8670 ;
      RECT 2.9230 0.8670 3.0530 0.9170 ;
      RECT 3.4310 0.5130 4.2970 0.5630 ;
      RECT 3.4310 0.5630 3.4810 0.6270 ;
      RECT 3.2270 0.6270 3.4810 0.6770 ;
      RECT 3.4310 0.6770 3.4810 1.0670 ;
      RECT 3.4310 1.0670 4.2970 1.1170 ;
      RECT 3.5310 0.6130 4.4330 0.6630 ;
      RECT 4.3830 0.3830 4.4330 0.6130 ;
      RECT 3.7350 0.6630 3.7850 0.9670 ;
      RECT 3.7350 0.9670 4.4330 1.0170 ;
      RECT 4.3830 1.0170 4.4330 1.2400 ;
      RECT 4.1390 0.7130 5.8930 0.7630 ;
      RECT 4.6870 0.7630 4.7370 1.2400 ;
      RECT 4.4950 0.5630 4.5450 0.7130 ;
      RECT 4.4950 0.5130 4.7370 0.5630 ;
      RECT 4.6870 0.3830 4.7370 0.5130 ;
      RECT 5.0670 0.6420 5.1170 0.7130 ;
      RECT 5.2190 0.6420 5.2690 0.7130 ;
      RECT 7.1190 0.4620 7.4130 0.5120 ;
      RECT 7.1190 0.1820 7.1690 0.4620 ;
      RECT 7.1190 0.5120 7.1690 0.6350 ;
      RECT 6.7990 0.1320 7.1690 0.1820 ;
      RECT 6.7990 0.6350 7.1690 0.6850 ;
      RECT 6.6630 0.4940 7.0170 0.5440 ;
      RECT 6.9670 0.3480 7.0170 0.4940 ;
      RECT 6.6630 0.5440 6.7130 0.7820 ;
      RECT 3.6830 1.5280 8.0230 1.5780 ;
      RECT 3.8350 0.7130 4.0690 0.7630 ;
      RECT 1.4790 0.9670 2.0930 1.0170 ;
      RECT 1.3430 0.4070 1.3930 0.6190 ;
      RECT 1.6470 0.6690 1.6970 0.9670 ;
      RECT 1.3430 0.6190 1.6970 0.6690 ;
      RECT 7.7270 0.5620 8.0210 0.6120 ;
      RECT 7.8620 0.4120 7.9120 0.5620 ;
      RECT 7.7270 0.3620 7.9120 0.4120 ;
      RECT 7.7270 0.6120 7.7770 0.8320 ;
      RECT 6.5630 0.8320 7.7770 0.8820 ;
      RECT 7.7270 0.1260 7.7770 0.3620 ;
      RECT 6.5630 0.4200 6.6130 0.8320 ;
      RECT 6.5630 0.3700 6.7310 0.4200 ;
      RECT 2.4670 0.8670 2.7210 0.9170 ;
      RECT 0.2790 0.6130 0.7250 0.6630 ;
      RECT 0.2790 0.8670 1.0290 0.9170 ;
      RECT 0.2790 0.4130 0.3290 0.6130 ;
      RECT 0.2790 0.6630 0.3290 0.8670 ;
      RECT 0.7190 0.5130 0.8610 0.5630 ;
      RECT 0.8110 0.5630 0.8610 0.6130 ;
      RECT 0.8110 0.6130 1.0290 0.6630 ;
      RECT 0.8110 0.6630 0.8610 0.7540 ;
      RECT 0.7180 0.7540 0.8610 0.8040 ;
      RECT 2.0110 0.6670 2.3970 0.7170 ;
      RECT 5.8110 1.2000 6.9570 1.2500 ;
      RECT 6.3590 1.0620 6.8050 1.1120 ;
      RECT 6.3590 0.1260 6.4090 1.0620 ;
  END
END RDFFNX2_LVT

MACRO RDFFSRARX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.208 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.4210 0.6630 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 8.2080 1.7020 ;
        RECT 0.2790 1.1310 0.3290 1.6420 ;
        RECT 0.8870 1.2940 0.9370 1.6420 ;
        RECT 2.1430 1.2700 2.1930 1.6420 ;
        RECT 6.2470 1.4540 6.2970 1.6420 ;
        RECT 0.7150 1.2440 0.9370 1.2940 ;
        RECT 1.9340 1.2200 3.0810 1.2700 ;
        RECT 3.7750 1.4040 6.2970 1.4540 ;
        RECT 3.7750 1.2790 3.8250 1.4040 ;
        RECT 4.8390 0.9590 4.8890 1.4040 ;
        RECT 4.3830 0.9530 4.4330 1.4040 ;
    END
  END VDD

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6870 0.4010 5.3870 0.4510 ;
        RECT 4.6870 0.1570 4.7370 0.4010 ;
        RECT 5.2650 0.4510 5.3870 0.5380 ;
        RECT 5.3370 0.5380 5.3870 0.8590 ;
        RECT 4.6870 0.8590 5.3870 0.9090 ;
        RECT 4.6870 0.9090 4.7370 1.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.9910 0.9690 5.5250 1.0190 ;
        RECT 5.4750 0.3510 5.5250 0.9690 ;
        RECT 4.9910 1.0190 5.2230 1.1290 ;
        RECT 4.9750 0.3010 5.5250 0.3510 ;
        RECT 4.9910 1.1290 5.0410 1.3270 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6430 1.4650 0.8150 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 8.2080 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.2720 ;
        RECT 4.8390 0.0300 4.8890 0.2410 ;
        RECT 6.8150 0.0300 6.8650 0.1980 ;
        RECT 7.2710 0.0300 7.3210 0.4260 ;
        RECT 5.9030 0.0300 5.9530 0.4260 ;
        RECT 4.5590 0.0300 4.6090 0.3000 ;
        RECT 0.2790 0.2720 2.1530 0.3220 ;
        RECT 3.7590 0.3000 4.6090 0.3500 ;
        RECT 1.9510 0.3220 2.0010 0.5570 ;
        RECT 0.7350 0.3220 0.7850 0.5570 ;
        RECT 0.8870 0.3220 0.9370 0.5570 ;
        RECT 2.1030 0.3220 2.1530 0.3280 ;
        RECT 0.2790 0.3220 0.3290 0.4050 ;
        RECT 2.1030 0.2440 2.1530 0.2720 ;
        RECT 2.1030 0.1940 3.0810 0.2440 ;
        RECT 2.4070 0.2440 2.4570 0.3490 ;
    END
  END VSS

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.2880 0.0930 4.3770 0.1430 ;
        RECT 4.3070 0.1430 4.3570 0.2000 ;
        RECT 3.8150 0.2000 4.3570 0.2500 ;
        RECT 3.8150 0.1380 3.8650 0.2000 ;
        RECT 1.6150 0.0880 3.8650 0.1380 ;
        RECT 1.6150 0.1380 1.7730 0.2100 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.3920 0.2490 7.5050 0.3590 ;
        RECT 7.4040 0.3590 7.4540 0.5270 ;
        RECT 7.1790 0.5270 7.4540 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6810 0.7030 2.8370 0.7310 ;
        RECT 2.6810 0.7310 3.1410 0.7810 ;
        RECT 2.7870 0.5970 2.8370 0.7030 ;
        RECT 2.6810 0.7810 2.8370 0.8150 ;
        RECT 3.0910 0.7810 3.1410 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 5.8870 0.9420 7.5050 1.0020 ;
        RECT 7.3950 0.6900 7.5050 0.9420 ;
        RECT 7.2710 0.6270 7.3210 0.9420 ;
    END
  END VDDG
  OBS
    LAYER PO ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 2.7970 0.0660 2.8270 0.6910 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 1.8850 0.9390 1.9150 1.6060 ;
      RECT 5.2290 0.0670 5.2590 1.6050 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 3.1010 0.8390 3.1310 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 3.8610 0.0660 3.8910 0.6910 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 3.7090 0.0660 3.7390 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 1.2770 0.8400 1.3070 1.6060 ;
      RECT 3.8610 0.9390 3.8910 1.6060 ;
      RECT 3.5570 0.0660 3.5870 0.6370 ;
      RECT 1.2770 0.0660 1.3070 0.6370 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 1.8850 0.0660 1.9150 0.6910 ;
      RECT 3.1010 0.0660 3.1310 0.6910 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 2.7970 0.8920 2.8270 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
      RECT 3.5570 0.8390 3.5870 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
    LAYER NWELL ;
      RECT 5.5840 0.4910 7.5950 1.0830 ;
      RECT -0.1150 1.5430 8.3300 1.7730 ;
      RECT -0.1150 0.6790 5.1220 1.5430 ;
      RECT 8.0550 0.6790 8.3300 1.5430 ;
    LAYER M1 ;
      RECT 3.3190 0.9670 3.5370 1.0170 ;
      RECT 3.3190 0.4440 3.3690 0.9670 ;
      RECT 3.3190 1.0170 3.3690 1.1200 ;
      RECT 2.8470 0.3940 3.5210 0.4440 ;
      RECT 3.4710 0.4440 3.5210 0.5630 ;
      RECT 3.4710 0.2970 3.5210 0.3940 ;
      RECT 3.3190 1.1700 3.3690 1.2700 ;
      RECT 2.8470 1.1200 3.3690 1.1700 ;
      RECT 2.2970 0.8580 2.3970 0.9080 ;
      RECT 2.2970 0.9080 2.3470 0.9680 ;
      RECT 1.8590 0.9680 2.3470 1.0180 ;
      RECT 1.3430 0.8540 2.2450 0.9040 ;
      RECT 1.3430 0.9040 1.3930 1.0590 ;
      RECT 1.3430 0.6130 1.3930 0.8540 ;
      RECT 1.3430 1.0590 1.7130 1.1090 ;
      RECT 1.3430 0.5630 1.5450 0.6130 ;
      RECT 1.3430 1.1090 1.3930 1.3370 ;
      RECT 1.4950 0.4070 1.5450 0.5630 ;
      RECT 1.3430 0.4130 1.3930 0.5630 ;
      RECT 4.4590 0.6320 4.8130 0.6820 ;
      RECT 4.7630 0.5970 4.8130 0.6320 ;
      RECT 3.9940 0.4500 4.0440 0.7290 ;
      RECT 3.9940 0.7290 4.1810 0.7790 ;
      RECT 4.1310 0.7790 4.1810 1.1790 ;
      RECT 3.6240 1.1790 4.1810 1.2290 ;
      RECT 4.4590 0.4500 4.5090 0.6320 ;
      RECT 3.6230 0.4000 4.5090 0.4500 ;
      RECT 3.6230 0.4500 3.6730 0.5630 ;
      RECT 3.6230 0.2970 3.6730 0.4000 ;
      RECT 3.6240 1.2290 3.6740 1.3530 ;
      RECT 4.8630 0.6130 5.2850 0.6630 ;
      RECT 4.2310 0.8090 4.2810 1.3010 ;
      RECT 4.2310 0.6780 4.2810 0.7590 ;
      RECT 4.1390 0.6280 4.2810 0.6780 ;
      RECT 4.2310 0.5000 4.2810 0.6280 ;
      RECT 4.5350 0.8090 4.5850 1.3010 ;
      RECT 4.8630 0.6630 4.9130 0.7590 ;
      RECT 4.2310 0.7590 4.9130 0.8090 ;
      RECT 5.2030 1.1990 6.5010 1.2490 ;
      RECT 3.4710 0.8670 3.6130 0.9170 ;
      RECT 3.4710 0.6630 3.5210 0.8670 ;
      RECT 3.4710 0.6130 3.9170 0.6630 ;
      RECT 3.1710 0.1880 3.7650 0.2380 ;
      RECT 3.1710 0.2380 3.2210 0.2940 ;
      RECT 2.5300 0.2940 3.2210 0.3440 ;
      RECT 2.1230 0.4550 2.1730 0.6130 ;
      RECT 1.8590 0.6130 2.1730 0.6630 ;
      RECT 2.5300 0.3440 2.5800 0.4050 ;
      RECT 2.1230 0.4050 2.5800 0.4550 ;
      RECT 3.7820 0.9670 3.9170 1.0170 ;
      RECT 3.7820 0.9160 3.8320 0.9670 ;
      RECT 3.6830 0.8660 3.8320 0.9160 ;
      RECT 3.2070 0.5440 3.2570 1.0200 ;
      RECT 2.6950 0.5170 3.2570 0.5440 ;
      RECT 2.7110 1.0200 3.2570 1.0700 ;
      RECT 2.6950 0.4940 3.2560 0.5170 ;
      RECT 2.4470 0.7880 2.4970 1.1200 ;
      RECT 1.5500 0.7380 2.4990 0.7880 ;
      RECT 2.2550 0.5050 2.3050 0.7380 ;
      RECT 2.7110 1.0700 2.7610 1.1200 ;
      RECT 2.2340 1.1200 2.7610 1.1700 ;
      RECT 1.1910 0.8130 1.2810 0.8630 ;
      RECT 1.2310 0.4620 1.2810 0.8130 ;
      RECT 1.1910 0.8630 1.2410 1.0830 ;
      RECT 1.1750 0.4120 1.2810 0.4620 ;
      RECT 0.4310 1.0830 1.2410 1.1330 ;
      RECT 1.1910 1.1330 1.2410 1.3540 ;
      RECT 0.4310 0.7980 0.4810 1.0830 ;
      RECT 0.4310 0.7480 0.5210 0.7980 ;
      RECT 0.4310 0.4350 0.5210 0.4850 ;
      RECT 0.4310 0.3720 0.4810 0.4350 ;
      RECT 0.4710 0.4850 0.5210 0.7480 ;
      RECT 0.5830 0.6130 1.0290 0.6630 ;
      RECT 0.5830 0.6630 0.6330 1.0040 ;
      RECT 0.5830 0.4130 0.6330 0.6130 ;
      RECT 0.7940 0.0940 1.4910 0.1440 ;
      RECT 6.1910 0.8200 6.7390 0.8700 ;
      RECT 6.4950 0.7090 7.0330 0.7590 ;
      RECT 7.1190 0.6770 7.1690 0.7680 ;
      RECT 7.0790 0.4270 7.1690 0.4620 ;
      RECT 7.1190 0.1260 7.1690 0.4270 ;
      RECT 7.0790 0.6270 7.1690 0.6770 ;
      RECT 7.0790 0.5120 7.1290 0.6270 ;
      RECT 6.8750 0.4770 7.1290 0.5120 ;
      RECT 6.8750 0.4620 7.1690 0.4770 ;
      RECT 6.4950 0.1320 6.7290 0.1820 ;
      RECT 5.7510 1.0620 6.2000 1.1120 ;
      RECT 5.7510 0.6770 5.8010 1.0620 ;
      RECT 5.7110 0.6270 5.8010 0.6770 ;
      RECT 5.7110 0.4770 5.7610 0.6270 ;
      RECT 5.7110 0.4270 5.8010 0.4770 ;
      RECT 5.7510 0.1260 5.8010 0.4270 ;
      RECT 1.0990 1.5240 2.0930 1.5740 ;
      RECT 5.8110 0.5270 6.4090 0.5770 ;
      RECT 6.0550 0.5770 6.1050 0.8840 ;
      RECT 6.0550 0.1260 6.1050 0.5270 ;
      RECT 6.3590 0.5770 6.4090 0.7700 ;
      RECT 6.3590 0.3480 6.4090 0.5270 ;
      RECT 3.9870 0.0940 4.2210 0.1440 ;
      RECT 6.7230 1.0570 7.2610 1.1070 ;
      RECT 6.1910 0.2480 7.0330 0.2980 ;
      RECT 3.2250 1.5200 6.1970 1.5700 ;
      RECT 2.4670 1.5200 3.1570 1.5700 ;
      RECT 2.9220 0.6130 3.1570 0.6630 ;
      RECT 2.5590 0.9200 2.9890 0.9700 ;
      RECT 2.9390 0.8310 2.9890 0.9200 ;
      RECT 2.5590 0.9700 2.6090 1.0340 ;
      RECT 2.5590 0.5050 2.6090 0.9200 ;
      RECT 2.3150 1.4200 3.6210 1.4700 ;
      RECT 1.4790 1.1900 1.8650 1.2400 ;
      RECT 1.4030 1.3890 1.9410 1.4390 ;
      RECT 1.0390 0.7130 1.1650 0.7630 ;
      RECT 1.0390 0.7630 1.0890 1.0330 ;
      RECT 1.1150 0.5630 1.1650 0.7130 ;
      RECT 1.0230 0.5130 1.1650 0.5630 ;
  END
END RDFFSRARX1_LVT

MACRO RDFFSRARX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.512 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.4210 0.6630 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 8.5120 1.7020 ;
        RECT 0.2790 1.1310 0.3290 1.6420 ;
        RECT 0.8870 1.2940 0.9370 1.6420 ;
        RECT 2.1430 1.2700 2.1930 1.6420 ;
        RECT 6.5510 1.4540 6.6010 1.6420 ;
        RECT 0.7150 1.2440 0.9370 1.2940 ;
        RECT 1.9340 1.2200 3.0810 1.2700 ;
        RECT 3.7750 1.4040 6.6010 1.4540 ;
        RECT 3.7750 1.2790 3.8250 1.4040 ;
        RECT 4.6870 0.9130 4.7370 1.4040 ;
        RECT 4.9910 0.9610 5.0410 1.4040 ;
        RECT 5.2950 1.0530 5.3450 1.4040 ;
        RECT 4.3830 0.9530 4.4330 1.4040 ;
    END
  END VDD

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6430 1.4650 0.8150 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 8.5120 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.2720 ;
        RECT 4.9910 0.0300 5.0410 0.3200 ;
        RECT 4.6870 0.0300 4.7370 0.4090 ;
        RECT 7.1190 0.0300 7.1690 0.1980 ;
        RECT 5.2950 0.0300 5.3450 0.2210 ;
        RECT 7.5750 0.0300 7.6250 0.4260 ;
        RECT 6.2070 0.0300 6.2570 0.4260 ;
        RECT 4.5590 0.0300 4.6090 0.3000 ;
        RECT 0.2790 0.2720 2.1530 0.3220 ;
        RECT 3.7590 0.3000 4.6090 0.3500 ;
        RECT 1.9510 0.3220 2.0010 0.5570 ;
        RECT 0.7350 0.3220 0.7850 0.5570 ;
        RECT 0.8870 0.3220 0.9370 0.5570 ;
        RECT 2.1030 0.3220 2.1530 0.3470 ;
        RECT 0.2790 0.3220 0.3290 0.4050 ;
        RECT 2.1030 0.2380 2.1530 0.2720 ;
        RECT 2.1030 0.1880 3.0810 0.2380 ;
        RECT 2.4070 0.2380 2.4570 0.3490 ;
    END
  END VSS

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6150 0.0970 3.8650 0.1380 ;
        RECT 1.6150 0.1380 1.7730 0.2100 ;
        RECT 3.8150 0.1380 3.8650 0.2000 ;
        RECT 1.7230 0.0880 3.8650 0.0970 ;
        RECT 3.8150 0.2000 4.3570 0.2500 ;
        RECT 4.3070 0.0880 4.3570 0.2000 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.5690 0.4000 5.6810 0.4020 ;
        RECT 4.8390 0.4020 5.6910 0.4520 ;
        RECT 4.8390 0.1490 4.8890 0.4020 ;
        RECT 5.5690 0.4520 5.6910 0.5120 ;
        RECT 5.6410 0.5120 5.6910 0.8420 ;
        RECT 4.8390 0.8420 5.6910 0.8920 ;
        RECT 4.8390 0.8920 4.8890 1.3190 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.6960 0.2490 7.8090 0.3590 ;
        RECT 7.7080 0.3590 7.7580 0.5270 ;
        RECT 7.4830 0.5270 7.7580 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6810 0.7050 2.8370 0.7310 ;
        RECT 2.6810 0.7310 3.1410 0.7810 ;
        RECT 2.7870 0.5970 2.8370 0.7050 ;
        RECT 2.6810 0.7810 2.8370 0.8150 ;
        RECT 3.0910 0.7810 3.1410 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 6.1910 0.9420 7.8090 1.0020 ;
        RECT 7.6990 0.6900 7.8090 0.9420 ;
        RECT 7.5750 0.6270 7.6250 0.9420 ;
    END
  END VDDG

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.1430 0.1490 5.1930 0.2710 ;
        RECT 5.1430 0.2710 5.8410 0.3210 ;
        RECT 5.7210 0.3210 5.8410 0.3600 ;
        RECT 5.7210 0.2500 5.8410 0.2710 ;
        RECT 5.7910 0.3600 5.8410 0.9420 ;
        RECT 5.7210 0.2470 5.8330 0.2500 ;
        RECT 5.1430 0.9420 5.8410 0.9920 ;
        RECT 5.1430 0.9920 5.1930 1.3270 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q
  OBS
    LAYER PO ;
      RECT 2.7970 0.0660 2.8270 0.6910 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 1.8850 0.9390 1.9150 1.6060 ;
      RECT 5.5330 0.0670 5.5630 1.6050 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 3.1010 0.8390 3.1310 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 3.8610 0.0660 3.8910 0.6910 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 3.7090 0.0660 3.7390 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 1.2770 0.8400 1.3070 1.6060 ;
      RECT 3.8610 0.9390 3.8910 1.6060 ;
      RECT 3.5570 0.0660 3.5870 0.6370 ;
      RECT 1.2770 0.0660 1.3070 0.6370 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 1.8850 0.0660 1.9150 0.6910 ;
      RECT 3.1010 0.0660 3.1310 0.6910 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 2.7970 0.8920 2.8270 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 3.5570 0.8390 3.5870 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
    LAYER NWELL ;
      RECT 5.8880 0.4910 7.8990 1.0830 ;
      RECT -0.1150 1.5430 8.6340 1.7730 ;
      RECT -0.1150 0.6790 5.4260 1.5430 ;
      RECT 8.3590 0.6790 8.6340 1.5430 ;
    LAYER M1 ;
      RECT 1.0390 0.7130 1.1650 0.7630 ;
      RECT 1.0390 0.7630 1.0890 1.0330 ;
      RECT 1.1150 0.5630 1.1650 0.7130 ;
      RECT 1.0230 0.5130 1.1650 0.5630 ;
      RECT 2.8470 0.3880 3.5210 0.4380 ;
      RECT 3.4710 0.4380 3.5210 0.5630 ;
      RECT 3.4710 0.2970 3.5210 0.3880 ;
      RECT 3.3190 0.4380 3.3690 0.9670 ;
      RECT 3.3190 0.9670 3.5370 1.0170 ;
      RECT 3.3190 1.0170 3.3690 1.1200 ;
      RECT 3.3190 1.1700 3.3690 1.2700 ;
      RECT 2.8470 1.1200 3.3690 1.1700 ;
      RECT 2.2970 0.8580 2.3970 0.9080 ;
      RECT 2.2970 0.9080 2.3470 0.9680 ;
      RECT 1.8590 0.9680 2.3470 1.0180 ;
      RECT 1.3430 0.8540 2.2450 0.9040 ;
      RECT 1.3430 0.9040 1.3930 1.0590 ;
      RECT 1.3430 0.6130 1.3930 0.8540 ;
      RECT 1.3430 1.0590 1.7130 1.1090 ;
      RECT 1.3430 0.5630 1.5450 0.6130 ;
      RECT 1.3430 1.1090 1.3930 1.3370 ;
      RECT 1.4950 0.4070 1.5450 0.5630 ;
      RECT 1.3430 0.4130 1.3930 0.5630 ;
      RECT 4.4590 0.6420 4.9810 0.6920 ;
      RECT 3.9940 0.4500 4.0440 0.7290 ;
      RECT 3.9940 0.7290 4.1810 0.7790 ;
      RECT 4.1310 0.7790 4.1810 1.1790 ;
      RECT 3.6240 1.1790 4.1810 1.2290 ;
      RECT 4.4590 0.4500 4.5090 0.6420 ;
      RECT 3.6230 0.4000 4.5090 0.4500 ;
      RECT 3.6230 0.4500 3.6730 0.5630 ;
      RECT 3.6230 0.2970 3.6730 0.4000 ;
      RECT 3.6240 1.2290 3.6740 1.3530 ;
      RECT 2.5590 0.9200 2.9890 0.9700 ;
      RECT 2.9390 0.8310 2.9890 0.9200 ;
      RECT 2.5590 0.9700 2.6090 1.0340 ;
      RECT 2.5590 0.5050 2.6090 0.9200 ;
      RECT 2.3150 1.4200 3.6210 1.4700 ;
      RECT 1.4790 1.1900 1.8650 1.2400 ;
      RECT 1.4030 1.3890 1.9410 1.4390 ;
      RECT 3.1710 0.1880 3.7650 0.2380 ;
      RECT 3.1710 0.2380 3.2210 0.2880 ;
      RECT 2.5300 0.2880 3.2210 0.3380 ;
      RECT 2.1230 0.4550 2.1730 0.6130 ;
      RECT 1.8590 0.6130 2.1730 0.6630 ;
      RECT 2.5300 0.3380 2.5800 0.4050 ;
      RECT 2.1230 0.4050 2.5800 0.4550 ;
      RECT 1.1910 0.8130 1.2810 0.8630 ;
      RECT 1.1910 0.8630 1.2410 1.0830 ;
      RECT 1.2310 0.4620 1.2810 0.8130 ;
      RECT 0.4310 1.0830 1.2410 1.1330 ;
      RECT 1.1750 0.4120 1.2810 0.4620 ;
      RECT 1.1910 1.1330 1.2410 1.3540 ;
      RECT 0.4310 0.7980 0.4810 1.0830 ;
      RECT 0.4310 0.7480 0.5210 0.7980 ;
      RECT 0.4310 0.4350 0.5210 0.4850 ;
      RECT 0.4310 0.3720 0.4810 0.4350 ;
      RECT 0.4710 0.4850 0.5210 0.7480 ;
      RECT 5.0310 0.6130 5.5890 0.6630 ;
      RECT 4.2310 0.7920 4.2810 1.3010 ;
      RECT 4.2310 0.6780 4.2810 0.7420 ;
      RECT 4.1390 0.6280 4.2810 0.6780 ;
      RECT 4.2310 0.5000 4.2810 0.6280 ;
      RECT 4.5350 0.7920 4.5850 1.3010 ;
      RECT 5.0310 0.6630 5.0810 0.7420 ;
      RECT 4.2310 0.7420 5.0810 0.7920 ;
      RECT 5.5070 1.1990 6.8050 1.2490 ;
      RECT 3.4710 0.8670 3.6130 0.9170 ;
      RECT 3.4710 0.6630 3.5210 0.8670 ;
      RECT 3.4710 0.6130 3.9170 0.6630 ;
      RECT 3.7820 0.9670 3.9170 1.0170 ;
      RECT 3.7820 0.9160 3.8320 0.9670 ;
      RECT 3.6830 0.8660 3.8320 0.9160 ;
      RECT 2.6950 0.4880 3.2570 0.5380 ;
      RECT 3.2070 0.5380 3.2570 1.0200 ;
      RECT 2.7110 1.0200 3.2570 1.0700 ;
      RECT 2.4470 0.7880 2.4970 1.1200 ;
      RECT 1.5500 0.7380 2.4990 0.7880 ;
      RECT 2.2550 0.5050 2.3050 0.7380 ;
      RECT 2.7110 1.0700 2.7610 1.1200 ;
      RECT 2.2340 1.1200 2.7610 1.1700 ;
      RECT 0.5830 0.6130 1.0290 0.6630 ;
      RECT 0.5830 0.6630 0.6330 1.0040 ;
      RECT 0.5830 0.4130 0.6330 0.6130 ;
      RECT 0.7940 0.0940 1.4910 0.1440 ;
      RECT 6.4950 0.8200 7.0430 0.8700 ;
      RECT 6.7990 0.7090 7.3370 0.7590 ;
      RECT 7.4230 0.6770 7.4730 0.7680 ;
      RECT 7.3830 0.4270 7.4730 0.4620 ;
      RECT 7.4230 0.1260 7.4730 0.4270 ;
      RECT 7.3830 0.6270 7.4730 0.6770 ;
      RECT 7.3830 0.5120 7.4330 0.6270 ;
      RECT 7.1790 0.4770 7.4330 0.5120 ;
      RECT 7.1790 0.4620 7.4730 0.4770 ;
      RECT 6.7990 0.1320 7.0330 0.1820 ;
      RECT 6.0550 1.0620 6.5040 1.1120 ;
      RECT 6.0550 0.6770 6.1050 1.0620 ;
      RECT 6.0150 0.6270 6.1050 0.6770 ;
      RECT 6.0150 0.4770 6.0650 0.6270 ;
      RECT 6.0150 0.4270 6.1050 0.4770 ;
      RECT 6.0550 0.1260 6.1050 0.4270 ;
      RECT 1.0990 1.5240 2.0930 1.5740 ;
      RECT 6.1150 0.5270 6.7130 0.5770 ;
      RECT 6.3590 0.5770 6.4090 0.8840 ;
      RECT 6.3590 0.1260 6.4090 0.5270 ;
      RECT 6.6630 0.5770 6.7130 0.7700 ;
      RECT 6.6630 0.3480 6.7130 0.5270 ;
      RECT 3.9870 0.0940 4.2210 0.1440 ;
      RECT 7.0270 1.0620 7.5650 1.1120 ;
      RECT 6.4950 0.2480 7.3370 0.2980 ;
      RECT 3.2250 1.5200 6.5010 1.5700 ;
      RECT 2.4670 1.5200 3.1570 1.5700 ;
      RECT 2.9220 0.6130 3.1570 0.6630 ;
  END
END RDFFSRARX2_LVT

MACRO RDFFSRASRX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.512 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 8.5120 1.7020 ;
        RECT 0.2790 1.1310 0.3290 1.6420 ;
        RECT 0.8870 1.2940 0.9370 1.6420 ;
        RECT 2.1430 1.2700 2.1930 1.6420 ;
        RECT 6.5510 1.4540 6.6010 1.6420 ;
        RECT 0.7150 1.2440 0.9370 1.2940 ;
        RECT 1.9340 1.2200 3.2330 1.2700 ;
        RECT 3.9270 1.4040 6.6010 1.4540 ;
        RECT 3.9270 1.2790 3.9770 1.4040 ;
        RECT 5.1430 1.0060 5.1930 1.4040 ;
        RECT 4.6870 0.9530 4.7370 1.4040 ;
    END
  END VDD

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.9910 0.4010 5.6910 0.4510 ;
        RECT 4.9910 0.1570 5.0410 0.4010 ;
        RECT 5.5690 0.4510 5.6910 0.5380 ;
        RECT 5.6410 0.5380 5.6910 0.8690 ;
        RECT 4.9910 0.8690 5.6910 0.9190 ;
        RECT 4.9910 0.9190 5.0410 1.3190 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2950 0.9790 5.8290 1.0290 ;
        RECT 5.2950 1.0290 5.5270 1.1290 ;
        RECT 5.7790 0.3510 5.8290 0.9790 ;
        RECT 5.2950 1.1290 5.3450 1.3370 ;
        RECT 5.2790 0.3010 5.8290 0.3510 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6430 1.4650 0.8150 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 8.5120 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.2640 ;
        RECT 5.1430 0.0300 5.1930 0.2410 ;
        RECT 7.1190 0.0300 7.1690 0.1980 ;
        RECT 7.5750 0.0300 7.6250 0.4260 ;
        RECT 6.2070 0.0300 6.2570 0.4260 ;
        RECT 4.8630 0.0300 4.9130 0.3000 ;
        RECT 0.2790 0.2640 2.1530 0.3140 ;
        RECT 3.9110 0.3000 4.9130 0.3500 ;
        RECT 1.9510 0.3140 2.0010 0.5570 ;
        RECT 0.7350 0.3140 0.7850 0.5570 ;
        RECT 0.8870 0.3140 0.9370 0.5570 ;
        RECT 2.1030 0.3140 2.1530 0.5330 ;
        RECT 0.2790 0.3140 0.3290 0.4050 ;
        RECT 2.1030 0.2470 2.1530 0.2640 ;
        RECT 2.1030 0.1970 3.2330 0.2470 ;
        RECT 2.5590 0.2470 2.6090 0.3490 ;
    END
  END VSS

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.1550 0.8570 4.3110 0.9750 ;
        RECT 4.1550 0.9750 4.2050 1.0790 ;
        RECT 3.6230 1.0790 4.2050 1.1290 ;
        RECT 3.6230 1.1290 3.6730 1.3200 ;
        RECT 2.3310 1.3200 3.6730 1.3700 ;
        RECT 2.3310 1.3700 2.3810 1.4550 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6150 0.0880 4.6610 0.1380 ;
        RECT 1.6150 0.1380 1.7730 0.2070 ;
        RECT 4.6110 0.1380 4.6610 0.1700 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.4210 0.6630 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.6970 0.2490 7.8090 0.3590 ;
        RECT 7.7080 0.3590 7.7580 0.5000 ;
        RECT 7.4830 0.5000 7.7580 0.5500 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8330 0.7050 2.9890 0.7310 ;
        RECT 2.8330 0.7310 3.2930 0.7810 ;
        RECT 2.9390 0.5970 2.9890 0.7050 ;
        RECT 2.8330 0.7810 2.9890 0.8150 ;
        RECT 3.2430 0.7810 3.2930 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 6.1910 0.9420 7.8090 1.0020 ;
        RECT 7.6990 0.6900 7.8090 0.9420 ;
        RECT 7.5750 0.6270 7.6250 0.9420 ;
    END
  END VDDG
  OBS
    LAYER PO ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 2.9490 0.0660 2.9790 0.6910 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 1.8850 0.9390 1.9150 1.6060 ;
      RECT 5.5330 0.0670 5.5630 1.6050 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 3.2530 0.8390 3.2830 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 4.0130 0.0660 4.0430 0.7360 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 1.2770 0.8400 1.3070 1.6060 ;
      RECT 4.0130 0.9390 4.0430 1.6060 ;
      RECT 3.7090 0.0660 3.7390 0.6530 ;
      RECT 1.2770 0.0660 1.3070 0.6370 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 1.8850 0.0660 1.9150 0.6910 ;
      RECT 3.2530 0.0660 3.2830 0.6910 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 2.9490 0.8920 2.9790 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 3.7090 0.8390 3.7390 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
    LAYER NWELL ;
      RECT 5.8880 0.4910 7.8990 1.0830 ;
      RECT -0.1150 1.5430 8.6340 1.7730 ;
      RECT -0.1150 0.6790 5.4260 1.5430 ;
      RECT 8.3590 0.6790 8.6340 1.5430 ;
    LAYER M1 ;
      RECT 1.0390 0.7130 1.1650 0.7630 ;
      RECT 1.0390 0.7630 1.0890 1.0330 ;
      RECT 1.1150 0.5630 1.1650 0.7130 ;
      RECT 1.0230 0.5130 1.1650 0.5630 ;
      RECT 2.9990 0.3970 3.6730 0.4470 ;
      RECT 3.6230 0.4470 3.6730 0.5630 ;
      RECT 3.6230 0.2970 3.6730 0.3970 ;
      RECT 3.4710 0.9670 3.6890 1.0170 ;
      RECT 3.4710 0.4470 3.5210 0.9670 ;
      RECT 3.4710 1.0170 3.5210 1.1200 ;
      RECT 3.4710 1.1700 3.5210 1.2700 ;
      RECT 2.9990 1.1200 3.5210 1.1700 ;
      RECT 2.3890 0.8580 2.5490 0.9080 ;
      RECT 2.3890 0.9080 2.4390 0.9680 ;
      RECT 1.8590 0.9680 2.4390 1.0180 ;
      RECT 1.3430 0.8540 2.2450 0.9040 ;
      RECT 1.3430 0.9040 1.3930 1.0590 ;
      RECT 1.3430 0.6130 1.3930 0.8540 ;
      RECT 1.3430 1.0590 1.7130 1.1090 ;
      RECT 1.3430 0.5630 1.5450 0.6130 ;
      RECT 1.3430 1.1090 1.3930 1.3370 ;
      RECT 1.4950 0.4070 1.5450 0.5630 ;
      RECT 1.3430 0.4130 1.3930 0.5630 ;
      RECT 4.7630 0.6690 5.1170 0.7190 ;
      RECT 5.0670 0.6340 5.1170 0.6690 ;
      RECT 4.1190 0.4500 4.1690 0.7570 ;
      RECT 4.4350 0.8070 4.4850 1.1790 ;
      RECT 4.7630 0.4500 4.8130 0.6690 ;
      RECT 3.7750 0.4000 4.8130 0.4500 ;
      RECT 3.7760 1.1790 4.4850 1.2290 ;
      RECT 4.1190 0.7570 4.4850 0.8070 ;
      RECT 3.7750 0.4500 3.8250 0.5630 ;
      RECT 3.7750 0.2970 3.8250 0.4000 ;
      RECT 3.7760 1.2290 3.8260 1.3530 ;
      RECT 1.1910 0.8130 1.2810 0.8630 ;
      RECT 1.1910 0.8630 1.2410 1.0830 ;
      RECT 1.2310 0.4620 1.2810 0.8130 ;
      RECT 0.4310 1.0830 1.2410 1.1330 ;
      RECT 1.1750 0.4120 1.2810 0.4620 ;
      RECT 1.1910 1.1330 1.2410 1.3540 ;
      RECT 0.4310 0.7980 0.4810 1.0830 ;
      RECT 0.4310 0.7480 0.5210 0.7980 ;
      RECT 0.4310 0.4350 0.5210 0.4850 ;
      RECT 0.4310 0.3720 0.4810 0.4350 ;
      RECT 0.4710 0.4850 0.5210 0.7480 ;
      RECT 3.3230 0.1970 3.9170 0.2470 ;
      RECT 3.3230 0.2470 3.3730 0.2970 ;
      RECT 2.6820 0.2970 3.3730 0.3470 ;
      RECT 2.2950 0.4550 2.3450 0.6130 ;
      RECT 1.8590 0.6130 2.3450 0.6630 ;
      RECT 2.6820 0.3470 2.7320 0.4050 ;
      RECT 2.2950 0.4050 2.7320 0.4550 ;
      RECT 5.1670 0.6130 5.5890 0.6630 ;
      RECT 4.5350 0.8190 4.5850 1.3010 ;
      RECT 4.5350 0.5500 4.5850 0.7690 ;
      RECT 4.3070 0.5000 4.5850 0.5500 ;
      RECT 4.3070 0.5500 4.3570 0.7070 ;
      RECT 4.8390 0.8190 4.8890 1.3010 ;
      RECT 5.1670 0.6630 5.2170 0.7690 ;
      RECT 4.5350 0.7690 5.2170 0.8190 ;
      RECT 5.5070 1.1990 6.8050 1.2490 ;
      RECT 3.6230 0.8670 3.7650 0.9170 ;
      RECT 3.6230 0.7040 3.6730 0.8670 ;
      RECT 3.6230 0.6540 4.0690 0.7040 ;
      RECT 3.9340 0.9670 4.0690 1.0170 ;
      RECT 3.9340 0.9160 3.9840 0.9670 ;
      RECT 3.8350 0.8660 3.9840 0.9160 ;
      RECT 2.8470 0.4970 3.4080 0.5070 ;
      RECT 3.3590 0.5470 3.4090 1.0200 ;
      RECT 2.8630 1.0200 3.4090 1.0700 ;
      RECT 2.8470 0.5070 3.4090 0.5470 ;
      RECT 2.5990 0.7880 2.6490 1.1200 ;
      RECT 1.5500 0.7380 2.6510 0.7880 ;
      RECT 2.4070 0.5050 2.4570 0.7380 ;
      RECT 2.8630 1.0700 2.9130 1.1200 ;
      RECT 2.0870 1.1200 2.9130 1.1700 ;
      RECT 0.5830 0.6130 1.0290 0.6630 ;
      RECT 0.5830 0.6630 0.6330 1.0040 ;
      RECT 0.5830 0.4130 0.6330 0.6130 ;
      RECT 0.7940 0.0940 1.4910 0.1440 ;
      RECT 6.4950 0.8200 7.0430 0.8700 ;
      RECT 6.7990 0.7090 7.3370 0.7590 ;
      RECT 7.3830 0.6270 7.4730 0.6770 ;
      RECT 7.4230 0.6770 7.4730 0.7680 ;
      RECT 7.3830 0.3910 7.4730 0.4410 ;
      RECT 7.4230 0.1260 7.4730 0.3910 ;
      RECT 7.3830 0.5120 7.4330 0.6270 ;
      RECT 7.1790 0.4620 7.4330 0.5120 ;
      RECT 7.3830 0.4410 7.4330 0.4620 ;
      RECT 6.7990 0.1320 7.0330 0.1820 ;
      RECT 6.0550 1.0700 6.5040 1.1200 ;
      RECT 6.0550 0.6770 6.1050 1.0700 ;
      RECT 6.0150 0.6270 6.1050 0.6770 ;
      RECT 6.0150 0.4770 6.0650 0.6270 ;
      RECT 6.0150 0.4270 6.1050 0.4770 ;
      RECT 6.0550 0.1260 6.1050 0.4270 ;
      RECT 1.0990 1.5240 2.0930 1.5740 ;
      RECT 6.1150 0.5270 6.7130 0.5770 ;
      RECT 6.3590 0.5770 6.4090 0.8690 ;
      RECT 6.3590 0.1260 6.4090 0.5270 ;
      RECT 6.6630 0.5770 6.7130 0.7700 ;
      RECT 6.6630 0.3480 6.7130 0.5270 ;
      RECT 7.0270 1.0910 7.5650 1.1410 ;
      RECT 6.4950 0.2480 7.3370 0.2980 ;
      RECT 3.3770 1.5200 6.5010 1.5700 ;
      RECT 2.6190 1.5200 3.3090 1.5700 ;
      RECT 3.0740 0.6130 3.3090 0.6630 ;
      RECT 2.7110 0.9200 3.1410 0.9700 ;
      RECT 3.0910 0.8310 3.1410 0.9200 ;
      RECT 2.7110 0.9700 2.7610 1.0340 ;
      RECT 2.7110 0.5050 2.7610 0.9200 ;
      RECT 2.4670 1.4200 3.7730 1.4700 ;
      RECT 1.4790 1.1900 1.8650 1.2400 ;
      RECT 4.0560 1.2870 4.4490 1.3370 ;
      RECT 1.4030 1.3890 1.9410 1.4390 ;
  END
END RDFFSRASRX1_LVT

MACRO RDFFSRASRX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.816 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 8.8160 1.7020 ;
        RECT 0.2790 1.1310 0.3290 1.6420 ;
        RECT 0.8870 1.2940 0.9370 1.6420 ;
        RECT 2.1430 1.2700 2.1930 1.6420 ;
        RECT 6.8550 1.4540 6.9050 1.6420 ;
        RECT 0.7150 1.2440 0.9370 1.2940 ;
        RECT 1.9340 1.2200 3.2330 1.2700 ;
        RECT 3.9270 1.4040 6.9050 1.4540 ;
        RECT 3.9270 1.2790 3.9770 1.4040 ;
        RECT 4.9910 0.9130 5.0410 1.4040 ;
        RECT 5.5990 1.0530 5.6490 1.4040 ;
        RECT 4.6870 0.9530 4.7370 1.4040 ;
        RECT 5.2950 0.9610 5.3450 1.4040 ;
    END
  END VDD

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6430 1.4650 0.8150 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 8.8160 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.2640 ;
        RECT 5.2950 0.0300 5.3450 0.3200 ;
        RECT 4.9910 0.0300 5.0410 0.4090 ;
        RECT 7.4230 0.0300 7.4730 0.1980 ;
        RECT 5.5990 0.0300 5.6490 0.2210 ;
        RECT 7.8790 0.0300 7.9290 0.4260 ;
        RECT 6.5110 0.0300 6.5610 0.4260 ;
        RECT 4.8630 0.0300 4.9130 0.2880 ;
        RECT 0.2790 0.2640 2.1530 0.3140 ;
        RECT 3.9110 0.2880 4.9130 0.3380 ;
        RECT 1.9510 0.3140 2.0010 0.5570 ;
        RECT 0.7350 0.3140 0.7850 0.5570 ;
        RECT 0.8870 0.3140 0.9370 0.5570 ;
        RECT 2.1030 0.3140 2.1530 0.5330 ;
        RECT 0.2790 0.3140 0.3290 0.4050 ;
        RECT 2.1030 0.2380 2.1530 0.2640 ;
        RECT 2.1030 0.1880 3.2330 0.2380 ;
        RECT 2.5590 0.2380 2.6090 0.3490 ;
    END
  END VSS

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.1550 0.8570 4.3110 0.9750 ;
        RECT 4.1550 0.9750 4.2050 1.0790 ;
        RECT 3.6230 1.0790 4.2050 1.1290 ;
        RECT 3.6230 1.1290 3.6730 1.3200 ;
        RECT 2.3310 1.3200 3.6730 1.3700 ;
        RECT 2.3310 1.3700 2.3810 1.4550 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6150 0.0880 4.6610 0.1380 ;
        RECT 1.6150 0.1380 1.7730 0.2100 ;
        RECT 4.6110 0.1380 4.6610 0.1700 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4470 0.1490 5.4970 0.2710 ;
        RECT 5.4470 0.2710 6.1450 0.3210 ;
        RECT 6.0250 0.3210 6.1450 0.3600 ;
        RECT 6.0250 0.2500 6.1450 0.2710 ;
        RECT 6.0950 0.3600 6.1450 0.9330 ;
        RECT 6.0250 0.2490 6.1370 0.2500 ;
        RECT 5.4470 0.9330 6.1450 0.9830 ;
        RECT 5.4470 0.9830 5.4970 1.3270 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.4210 0.6630 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8730 0.4000 5.9850 0.4020 ;
        RECT 5.1430 0.4020 5.9950 0.4520 ;
        RECT 5.1430 0.1490 5.1930 0.4020 ;
        RECT 5.8730 0.4520 5.9950 0.5120 ;
        RECT 5.9450 0.5120 5.9950 0.8330 ;
        RECT 5.1430 0.8330 5.9950 0.8830 ;
        RECT 5.1430 0.8830 5.1930 1.3190 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.0010 0.2490 8.1130 0.3590 ;
        RECT 8.0120 0.3590 8.0620 0.5270 ;
        RECT 7.7870 0.5270 8.0620 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8330 0.7050 2.9890 0.7310 ;
        RECT 2.8330 0.7310 3.2930 0.7810 ;
        RECT 2.9390 0.5970 2.9890 0.7050 ;
        RECT 2.8330 0.7810 2.9890 0.8150 ;
        RECT 3.2430 0.7810 3.2930 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 6.4950 0.9420 8.1130 1.0020 ;
        RECT 8.0030 0.6900 8.1130 0.9420 ;
        RECT 7.8790 0.6270 7.9290 0.9420 ;
    END
  END VDDG
  OBS
    LAYER PO ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 2.9490 0.0660 2.9790 0.6910 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 1.8850 0.9390 1.9150 1.6060 ;
      RECT 5.8370 0.0670 5.8670 1.6050 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 3.2530 0.8390 3.2830 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 4.0130 0.0660 4.0430 0.6910 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 1.2770 0.8400 1.3070 1.6060 ;
      RECT 4.0130 0.9390 4.0430 1.6060 ;
      RECT 3.7090 0.0660 3.7390 0.6370 ;
      RECT 1.2770 0.0660 1.3070 0.6370 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
      RECT 1.8850 0.0660 1.9150 0.6910 ;
      RECT 3.2530 0.0660 3.2830 0.6910 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 2.9490 0.8920 2.9790 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 3.7090 0.8390 3.7390 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
    LAYER NWELL ;
      RECT 6.1920 0.4910 8.2030 1.0830 ;
      RECT -0.1150 1.5430 8.9380 1.7730 ;
      RECT -0.1150 0.6790 5.7300 1.5430 ;
      RECT 8.6630 0.6790 8.9380 1.5430 ;
    LAYER M1 ;
      RECT 1.0390 0.7130 1.1650 0.7630 ;
      RECT 1.0390 0.7630 1.0890 1.0330 ;
      RECT 1.1150 0.5630 1.1650 0.7130 ;
      RECT 1.0230 0.5130 1.1650 0.5630 ;
      RECT 2.9990 0.3880 3.6730 0.4380 ;
      RECT 3.6230 0.4380 3.6730 0.5630 ;
      RECT 3.6230 0.2970 3.6730 0.3880 ;
      RECT 3.4710 0.9670 3.6890 1.0170 ;
      RECT 3.4710 0.4380 3.5210 0.9670 ;
      RECT 3.4710 1.0170 3.5210 1.1200 ;
      RECT 3.4710 1.1700 3.5210 1.2700 ;
      RECT 2.9990 1.1200 3.5210 1.1700 ;
      RECT 2.3890 0.8580 2.5490 0.9080 ;
      RECT 2.3890 0.9080 2.4390 0.9680 ;
      RECT 1.8590 0.9680 2.4390 1.0180 ;
      RECT 1.3430 0.8540 2.2450 0.9040 ;
      RECT 1.3430 0.9040 1.3930 1.0590 ;
      RECT 1.3430 0.6130 1.3930 0.8540 ;
      RECT 1.3430 1.0590 1.7130 1.1090 ;
      RECT 1.3430 0.5630 1.5450 0.6130 ;
      RECT 1.3430 1.1090 1.3930 1.3370 ;
      RECT 1.4950 0.4070 1.5450 0.5630 ;
      RECT 1.3430 0.4130 1.3930 0.5630 ;
      RECT 4.7320 0.6320 5.2850 0.6820 ;
      RECT 4.1190 0.4500 4.1690 0.7290 ;
      RECT 4.1190 0.7290 4.4850 0.7790 ;
      RECT 4.4350 0.7790 4.4850 1.1790 ;
      RECT 4.7630 0.4500 4.8130 0.6320 ;
      RECT 3.7750 0.4000 4.8130 0.4500 ;
      RECT 3.7760 1.1790 4.4850 1.2290 ;
      RECT 3.7750 0.4500 3.8250 0.5630 ;
      RECT 3.7750 0.2970 3.8250 0.4000 ;
      RECT 3.7760 1.2290 3.8260 1.3530 ;
      RECT 3.3590 0.5380 3.4090 1.0200 ;
      RECT 2.8470 0.5110 3.4090 0.5380 ;
      RECT 2.8630 1.0200 3.4090 1.0700 ;
      RECT 2.8470 0.4880 3.4080 0.5110 ;
      RECT 2.5990 0.7880 2.6490 1.1200 ;
      RECT 1.5500 0.7380 2.6510 0.7880 ;
      RECT 2.4070 0.5050 2.4570 0.7380 ;
      RECT 2.8630 1.0700 2.9130 1.1200 ;
      RECT 2.0870 1.1200 2.9130 1.1700 ;
      RECT 3.6230 0.8670 3.7650 0.9170 ;
      RECT 3.6230 0.6630 3.6730 0.8670 ;
      RECT 3.6230 0.6130 4.0690 0.6630 ;
      RECT 2.7110 0.9200 3.1410 0.9700 ;
      RECT 3.0910 0.8310 3.1410 0.9200 ;
      RECT 2.7110 0.9700 2.7610 1.0340 ;
      RECT 2.7110 0.5050 2.7610 0.9200 ;
      RECT 2.4670 1.4200 3.7730 1.4700 ;
      RECT 1.4790 1.1900 1.8650 1.2400 ;
      RECT 4.0560 1.2870 4.4490 1.3370 ;
      RECT 1.4030 1.3890 1.9410 1.4390 ;
      RECT 3.3230 0.1880 3.9170 0.2380 ;
      RECT 3.3230 0.2380 3.3730 0.2880 ;
      RECT 2.6820 0.2880 3.3730 0.3380 ;
      RECT 2.2950 0.4550 2.3450 0.6130 ;
      RECT 1.8590 0.6130 2.3450 0.6630 ;
      RECT 2.6820 0.3380 2.7320 0.4050 ;
      RECT 2.2950 0.4050 2.7320 0.4550 ;
      RECT 1.1910 0.8130 1.2810 0.8630 ;
      RECT 1.1910 0.8630 1.2410 1.0830 ;
      RECT 1.2310 0.4620 1.2810 0.8130 ;
      RECT 0.4310 1.0830 1.2410 1.1330 ;
      RECT 1.1750 0.4120 1.2810 0.4620 ;
      RECT 1.1910 1.1330 1.2410 1.3540 ;
      RECT 0.4310 0.7980 0.4810 1.0830 ;
      RECT 0.4310 0.7480 0.5210 0.7980 ;
      RECT 0.4310 0.4350 0.5210 0.4850 ;
      RECT 0.4310 0.3720 0.4810 0.4350 ;
      RECT 0.4710 0.4850 0.5210 0.7480 ;
      RECT 5.3440 0.6130 5.8930 0.6630 ;
      RECT 4.5350 0.7830 4.5850 1.3010 ;
      RECT 4.5350 0.5500 4.5850 0.7330 ;
      RECT 4.3070 0.5000 4.5850 0.5500 ;
      RECT 4.3070 0.5500 4.3570 0.6790 ;
      RECT 4.8390 0.7830 4.8890 1.3010 ;
      RECT 5.3440 0.6630 5.3940 0.7330 ;
      RECT 4.5350 0.7330 5.3940 0.7830 ;
      RECT 5.8110 1.1990 7.1090 1.2490 ;
      RECT 3.9340 0.9670 4.0690 1.0170 ;
      RECT 3.9340 0.9160 3.9840 0.9670 ;
      RECT 3.8350 0.8660 3.9840 0.9160 ;
      RECT 0.5830 0.6130 1.0290 0.6630 ;
      RECT 0.5830 0.6630 0.6330 1.0040 ;
      RECT 0.5830 0.4130 0.6330 0.6130 ;
      RECT 0.7940 0.0940 1.4910 0.1440 ;
      RECT 6.7990 0.8200 7.3470 0.8700 ;
      RECT 7.1030 0.7090 7.6410 0.7590 ;
      RECT 7.7270 0.6770 7.7770 0.7680 ;
      RECT 7.6870 0.4270 7.7770 0.4620 ;
      RECT 7.7270 0.1260 7.7770 0.4270 ;
      RECT 7.6870 0.6270 7.7770 0.6770 ;
      RECT 7.6870 0.5120 7.7370 0.6270 ;
      RECT 7.4830 0.4770 7.7370 0.5120 ;
      RECT 7.4830 0.4620 7.7770 0.4770 ;
      RECT 7.1030 0.1320 7.3370 0.1820 ;
      RECT 6.3590 1.0620 6.8080 1.1120 ;
      RECT 6.3590 0.6770 6.4090 1.0620 ;
      RECT 6.3190 0.6270 6.4090 0.6770 ;
      RECT 6.3190 0.4770 6.3690 0.6270 ;
      RECT 6.3190 0.4270 6.4090 0.4770 ;
      RECT 6.3590 0.1260 6.4090 0.4270 ;
      RECT 1.0990 1.5240 2.0930 1.5740 ;
      RECT 6.4190 0.5270 7.0170 0.5770 ;
      RECT 6.6630 0.5770 6.7130 0.8840 ;
      RECT 6.6630 0.1210 6.7130 0.5270 ;
      RECT 6.9670 0.5770 7.0170 0.7700 ;
      RECT 6.9670 0.3480 7.0170 0.5270 ;
      RECT 7.3310 1.0620 7.8690 1.1120 ;
      RECT 6.7990 0.2480 7.6410 0.2980 ;
      RECT 3.3770 1.5200 6.8050 1.5700 ;
      RECT 2.6190 1.5200 3.3090 1.5700 ;
      RECT 3.0740 0.6130 3.3090 0.6630 ;
  END
END RDFFSRASRX2_LVT

MACRO RDFFSRASX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.512 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 8.5120 1.7020 ;
        RECT 0.2790 1.1310 0.3290 1.6420 ;
        RECT 0.8870 1.2940 0.9370 1.6420 ;
        RECT 2.1430 1.2700 2.1930 1.6420 ;
        RECT 6.5510 1.4540 6.6010 1.6420 ;
        RECT 0.7150 1.2440 0.9370 1.2940 ;
        RECT 1.9340 1.2200 3.2330 1.2700 ;
        RECT 3.9270 1.4040 6.6010 1.4540 ;
        RECT 3.9270 1.2790 3.9770 1.4040 ;
        RECT 5.1430 0.9590 5.1930 1.4040 ;
        RECT 4.6870 0.9530 4.7370 1.4040 ;
    END
  END VDD

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.9910 0.4010 5.6910 0.4510 ;
        RECT 4.9910 0.1570 5.0410 0.4010 ;
        RECT 5.5690 0.4510 5.6910 0.5380 ;
        RECT 5.6410 0.5380 5.6910 0.8590 ;
        RECT 4.9910 0.8590 5.6910 0.9090 ;
        RECT 4.9910 0.9090 5.0410 1.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2950 0.9690 5.8290 1.0190 ;
        RECT 5.7790 0.3510 5.8290 0.9690 ;
        RECT 5.2950 1.0190 5.5270 1.1290 ;
        RECT 5.2790 0.3010 5.8290 0.3510 ;
        RECT 5.2950 1.1290 5.3450 1.3270 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6430 1.4650 0.8150 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 8.5120 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.2720 ;
        RECT 5.1430 0.0300 5.1930 0.2410 ;
        RECT 7.1190 0.0300 7.1690 0.1980 ;
        RECT 7.5750 0.0300 7.6250 0.4260 ;
        RECT 6.2070 0.0300 6.2570 0.4260 ;
        RECT 4.8630 0.0300 4.9130 0.2880 ;
        RECT 0.2790 0.2720 2.1530 0.3220 ;
        RECT 3.9110 0.2880 4.9130 0.3380 ;
        RECT 1.9510 0.3220 2.0010 0.5570 ;
        RECT 0.7350 0.3220 0.7850 0.5570 ;
        RECT 0.8870 0.3220 0.9370 0.5570 ;
        RECT 2.1030 0.3220 2.1530 0.5330 ;
        RECT 0.2790 0.3220 0.3290 0.4050 ;
        RECT 2.1030 0.2380 2.1530 0.2720 ;
        RECT 2.1030 0.1880 3.2330 0.2380 ;
        RECT 2.5590 0.2380 2.6090 0.3490 ;
    END
  END VSS

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.1550 0.8570 4.3110 0.9750 ;
        RECT 4.1550 0.9750 4.2050 1.0790 ;
        RECT 3.6230 1.0790 4.2050 1.1290 ;
        RECT 3.6230 1.1290 3.6730 1.3200 ;
        RECT 2.3310 1.3200 3.6730 1.3700 ;
        RECT 2.3310 1.3700 2.3810 1.4550 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.4210 0.6630 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.6970 0.2490 7.8090 0.3590 ;
        RECT 7.7080 0.3590 7.7580 0.5170 ;
        RECT 7.4830 0.5170 7.7580 0.5670 ;
        RECT 7.7080 0.5670 7.7580 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8330 0.7040 2.9890 0.7310 ;
        RECT 2.8330 0.7310 3.2930 0.7810 ;
        RECT 2.9390 0.5970 2.9890 0.7040 ;
        RECT 2.8330 0.7810 2.9890 0.8150 ;
        RECT 3.2430 0.7810 3.2930 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 6.1910 0.9420 7.8090 1.0020 ;
        RECT 7.6990 0.6900 7.8090 0.9420 ;
        RECT 7.5750 0.6270 7.6250 0.9420 ;
    END
  END VDDG
  OBS
    LAYER PO ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 2.9490 0.0660 2.9790 0.6910 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 1.8850 0.9390 1.9150 1.6060 ;
      RECT 5.5330 0.0670 5.5630 1.6050 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 3.2530 0.8390 3.2830 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 4.0130 0.0660 4.0430 0.6910 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 1.2770 0.8400 1.3070 1.6060 ;
      RECT 4.0130 0.9390 4.0430 1.6060 ;
      RECT 3.7090 0.0660 3.7390 0.6370 ;
      RECT 1.2770 0.0660 1.3070 0.6370 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 1.8850 0.0660 1.9150 0.6910 ;
      RECT 3.2530 0.0660 3.2830 0.6910 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 2.9490 0.8920 2.9790 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 3.7090 0.8390 3.7390 1.6060 ;
    LAYER NWELL ;
      RECT 5.8880 0.4910 7.8990 1.0830 ;
      RECT -0.1150 1.5430 8.6340 1.7730 ;
      RECT -0.1150 0.6790 5.4260 1.5430 ;
      RECT 8.3590 0.6790 8.6340 1.5430 ;
    LAYER M1 ;
      RECT 1.0390 0.7630 1.0890 1.0330 ;
      RECT 1.0390 0.7130 1.1650 0.7630 ;
      RECT 1.1150 0.5630 1.1650 0.7130 ;
      RECT 1.0230 0.5130 1.1650 0.5630 ;
      RECT 2.9990 0.3880 3.6730 0.4380 ;
      RECT 3.6230 0.4380 3.6730 0.5630 ;
      RECT 3.6230 0.2970 3.6730 0.3880 ;
      RECT 3.4710 0.9670 3.6890 1.0170 ;
      RECT 3.4710 0.3840 3.5210 0.3880 ;
      RECT 3.4710 0.4380 3.5210 0.9670 ;
      RECT 3.4710 1.0170 3.5210 1.1200 ;
      RECT 3.4710 1.1700 3.5210 1.2700 ;
      RECT 2.9990 1.1200 3.5210 1.1700 ;
      RECT 2.3890 0.8580 2.5490 0.9080 ;
      RECT 2.3890 0.9080 2.4390 0.9680 ;
      RECT 1.8590 0.9680 2.4390 1.0180 ;
      RECT 1.3430 0.8540 2.2450 0.9040 ;
      RECT 1.3430 0.9040 1.3930 1.0590 ;
      RECT 1.3430 0.6130 1.3930 0.8540 ;
      RECT 1.3430 1.0590 1.7130 1.1090 ;
      RECT 1.3430 0.5630 1.5450 0.6130 ;
      RECT 1.3430 1.1090 1.3930 1.3370 ;
      RECT 1.4950 0.4070 1.5450 0.5630 ;
      RECT 1.3430 0.4130 1.3930 0.5630 ;
      RECT 4.7630 0.6420 5.1170 0.6920 ;
      RECT 5.0670 0.5970 5.1170 0.6420 ;
      RECT 4.1190 0.4500 4.1690 0.7290 ;
      RECT 4.1190 0.7290 4.4850 0.7790 ;
      RECT 4.4350 0.7790 4.4850 1.1790 ;
      RECT 4.7630 0.4500 4.8130 0.6420 ;
      RECT 3.7750 0.4000 4.8130 0.4500 ;
      RECT 3.7760 1.1790 4.4850 1.2290 ;
      RECT 3.7750 0.4500 3.8250 0.5630 ;
      RECT 3.7750 0.2970 3.8250 0.4000 ;
      RECT 3.7760 1.2290 3.8260 1.3530 ;
      RECT 1.1910 0.8130 1.2810 0.8630 ;
      RECT 1.1910 0.8630 1.2410 1.0830 ;
      RECT 1.2310 0.4620 1.2810 0.8130 ;
      RECT 0.4310 1.0830 1.2410 1.1330 ;
      RECT 1.1750 0.4120 1.2810 0.4620 ;
      RECT 1.1910 1.1330 1.2410 1.3540 ;
      RECT 0.4310 0.7980 0.4810 1.0830 ;
      RECT 0.4310 0.7480 0.5210 0.7980 ;
      RECT 0.4310 0.4350 0.5210 0.4850 ;
      RECT 0.4310 0.3720 0.4810 0.4350 ;
      RECT 0.4710 0.4850 0.5210 0.7480 ;
      RECT 3.3230 0.1880 3.9170 0.2380 ;
      RECT 3.3230 0.2380 3.3730 0.2880 ;
      RECT 2.6820 0.2880 3.3730 0.3380 ;
      RECT 2.2950 0.4550 2.3450 0.6130 ;
      RECT 1.8590 0.6130 2.3450 0.6630 ;
      RECT 2.6820 0.3380 2.7320 0.4050 ;
      RECT 2.2950 0.4050 2.7320 0.4550 ;
      RECT 5.1670 0.6130 5.5890 0.6630 ;
      RECT 4.5350 0.8090 4.5850 1.3010 ;
      RECT 4.5350 0.5500 4.5850 0.7590 ;
      RECT 4.3070 0.5000 4.5850 0.5500 ;
      RECT 4.3070 0.5500 4.3570 0.6790 ;
      RECT 4.8390 0.8090 4.8890 1.3010 ;
      RECT 5.1670 0.6630 5.2170 0.7590 ;
      RECT 4.5350 0.7590 5.2170 0.8090 ;
      RECT 5.5070 1.1990 6.8050 1.2490 ;
      RECT 3.6230 0.8670 3.7650 0.9170 ;
      RECT 3.6230 0.6630 3.6730 0.8670 ;
      RECT 3.6230 0.6130 4.0690 0.6630 ;
      RECT 3.9340 0.9670 4.0690 1.0170 ;
      RECT 3.9340 0.9160 3.9840 0.9670 ;
      RECT 3.8350 0.8660 3.9840 0.9160 ;
      RECT 2.8470 0.4880 3.4080 0.5070 ;
      RECT 2.8470 0.5070 3.4090 0.5380 ;
      RECT 3.3590 0.5380 3.4090 1.0200 ;
      RECT 2.8630 1.0200 3.4090 1.0700 ;
      RECT 2.5990 0.7880 2.6490 1.1200 ;
      RECT 1.5500 0.7380 2.6510 0.7880 ;
      RECT 2.4070 0.5050 2.4570 0.7380 ;
      RECT 2.8630 1.0700 2.9130 1.1200 ;
      RECT 2.0870 1.1200 2.9130 1.1700 ;
      RECT 0.5830 0.6130 1.0290 0.6630 ;
      RECT 0.5830 0.6630 0.6330 1.0040 ;
      RECT 0.5830 0.4130 0.6330 0.6130 ;
      RECT 0.7940 0.0940 1.4910 0.1440 ;
      RECT 4.6110 0.1380 4.6610 0.1700 ;
      RECT 1.7230 0.0880 4.6610 0.1380 ;
      RECT 1.7230 0.1380 1.7730 0.1700 ;
      RECT 6.4950 0.8200 7.0430 0.8700 ;
      RECT 6.7990 0.7090 7.3370 0.7590 ;
      RECT 7.3830 0.6270 7.4730 0.6770 ;
      RECT 7.4230 0.6770 7.4730 0.7680 ;
      RECT 7.3830 0.4580 7.4330 0.4620 ;
      RECT 7.3830 0.4080 7.4730 0.4580 ;
      RECT 7.4230 0.1260 7.4730 0.4080 ;
      RECT 7.3830 0.5120 7.4330 0.6270 ;
      RECT 7.1790 0.4620 7.4330 0.5120 ;
      RECT 6.7990 0.1320 7.0330 0.1820 ;
      RECT 6.0550 1.0620 6.5040 1.1120 ;
      RECT 6.0550 0.6770 6.1050 1.0620 ;
      RECT 6.0150 0.6270 6.1050 0.6770 ;
      RECT 6.0150 0.4770 6.0650 0.6270 ;
      RECT 6.0150 0.4270 6.1050 0.4770 ;
      RECT 6.0550 0.1260 6.1050 0.4270 ;
      RECT 1.0990 1.5240 2.0930 1.5740 ;
      RECT 6.1150 0.5270 6.7130 0.5770 ;
      RECT 6.3590 0.5770 6.4090 0.8840 ;
      RECT 6.3590 0.1260 6.4090 0.5270 ;
      RECT 6.6630 0.5770 6.7130 0.7700 ;
      RECT 6.6630 0.3480 6.7130 0.5270 ;
      RECT 7.0270 1.0620 7.5650 1.1120 ;
      RECT 6.4950 0.2480 7.3370 0.2980 ;
      RECT 3.3770 1.5200 6.5010 1.5700 ;
      RECT 2.6190 1.5200 3.3090 1.5700 ;
      RECT 3.0740 0.6130 3.3090 0.6630 ;
      RECT 2.7110 0.9200 3.1410 0.9700 ;
      RECT 3.0910 0.8310 3.1410 0.9200 ;
      RECT 2.7110 0.9700 2.7610 1.0340 ;
      RECT 2.7110 0.5050 2.7610 0.9200 ;
      RECT 2.4670 1.4200 3.7730 1.4700 ;
      RECT 1.4790 1.1900 1.8650 1.2400 ;
      RECT 4.0560 1.2790 4.4490 1.3290 ;
      RECT 1.4030 1.3890 1.9410 1.4390 ;
  END
END RDFFSRASX1_LVT

MACRO RDFFSRASX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.816 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8730 0.4010 5.9850 0.4020 ;
        RECT 5.1430 0.4020 5.9950 0.4520 ;
        RECT 5.1430 0.1490 5.1930 0.4020 ;
        RECT 5.8730 0.4520 5.9950 0.5120 ;
        RECT 5.9450 0.5120 5.9950 0.8420 ;
        RECT 5.1430 0.8420 5.9950 0.8920 ;
        RECT 5.1430 0.8920 5.1930 1.3190 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4470 0.2710 6.1450 0.3210 ;
        RECT 6.0250 0.3210 6.1450 0.3600 ;
        RECT 6.0250 0.2500 6.1450 0.2710 ;
        RECT 5.4470 0.1490 5.4970 0.2710 ;
        RECT 6.0950 0.3600 6.1450 0.9420 ;
        RECT 6.0250 0.2490 6.1370 0.2500 ;
        RECT 5.4470 0.9420 6.1450 0.9920 ;
        RECT 5.4470 0.9920 5.4970 1.3270 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 8.8160 1.7020 ;
        RECT 0.2790 1.1310 0.3290 1.6420 ;
        RECT 0.8870 1.2940 0.9370 1.6420 ;
        RECT 2.1430 1.2700 2.1930 1.6420 ;
        RECT 6.8550 1.4540 6.9050 1.6420 ;
        RECT 0.7150 1.2440 0.9370 1.2940 ;
        RECT 1.9340 1.2200 3.2330 1.2700 ;
        RECT 3.9270 1.4040 6.9050 1.4540 ;
        RECT 3.9270 1.2790 3.9770 1.4040 ;
        RECT 4.6870 0.9530 4.7370 1.4040 ;
        RECT 5.2950 0.9610 5.3450 1.4040 ;
        RECT 4.9910 0.9130 5.0410 1.4040 ;
        RECT 5.5990 1.0530 5.6490 1.4040 ;
    END
  END VDD

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6430 1.4650 0.8150 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 8.8160 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.2720 ;
        RECT 5.2950 0.0300 5.3450 0.3200 ;
        RECT 4.9910 0.0300 5.0410 0.4090 ;
        RECT 5.5990 0.0300 5.6490 0.2210 ;
        RECT 6.5110 0.0300 6.5610 0.4260 ;
        RECT 7.4230 0.0300 7.4730 0.1980 ;
        RECT 7.8790 0.0300 7.9290 0.4260 ;
        RECT 4.8630 0.0300 4.9130 0.2880 ;
        RECT 0.2790 0.2720 2.1530 0.3220 ;
        RECT 3.9110 0.2880 4.9130 0.3380 ;
        RECT 1.9510 0.3220 2.0010 0.5570 ;
        RECT 0.7350 0.3220 0.7850 0.5570 ;
        RECT 0.8870 0.3220 0.9370 0.5570 ;
        RECT 2.1030 0.3220 2.1530 0.5330 ;
        RECT 0.2790 0.3220 0.3290 0.4050 ;
        RECT 2.1030 0.2380 2.1530 0.2720 ;
        RECT 2.1030 0.1880 3.2330 0.2380 ;
        RECT 2.5590 0.2380 2.6090 0.3490 ;
    END
  END VSS

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.1550 0.8570 4.3110 0.9750 ;
        RECT 4.1550 0.9750 4.2050 1.0790 ;
        RECT 3.6230 1.0790 4.2050 1.1290 ;
        RECT 3.6230 1.1290 3.6730 1.3200 ;
        RECT 2.3310 1.3200 3.6730 1.3700 ;
        RECT 2.3310 1.3700 2.3810 1.4550 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.4210 0.6630 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.0010 0.2490 8.1130 0.3590 ;
        RECT 8.0120 0.3590 8.0620 0.5270 ;
        RECT 7.7870 0.5270 8.0620 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8330 0.7050 2.9890 0.7310 ;
        RECT 2.8330 0.7310 3.2930 0.7810 ;
        RECT 2.9390 0.5970 2.9890 0.7050 ;
        RECT 2.8330 0.7810 2.9890 0.8150 ;
        RECT 3.2430 0.7810 3.2930 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 6.4950 0.9420 8.1130 1.0020 ;
        RECT 8.0030 0.6900 8.1130 0.9420 ;
        RECT 7.8790 0.6270 7.9290 0.9420 ;
    END
  END VDDG
  OBS
    LAYER PO ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 2.9490 0.0660 2.9790 0.6910 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 1.8850 0.9390 1.9150 1.6060 ;
      RECT 5.8370 0.0670 5.8670 1.6050 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 3.2530 0.8390 3.2830 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 4.0130 0.0660 4.0430 0.6910 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 1.2770 0.8400 1.3070 1.6060 ;
      RECT 4.0130 0.9390 4.0430 1.6060 ;
      RECT 3.7090 0.0660 3.7390 0.6370 ;
      RECT 1.2770 0.0660 1.3070 0.6370 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
      RECT 1.8850 0.0660 1.9150 0.6910 ;
      RECT 3.2530 0.0660 3.2830 0.6910 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 2.9490 0.8920 2.9790 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 3.7090 0.8390 3.7390 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
    LAYER NWELL ;
      RECT 6.1920 0.4910 8.2030 1.0830 ;
      RECT -0.1150 1.5430 8.9380 1.7730 ;
      RECT -0.1150 0.6790 5.7300 1.5430 ;
      RECT 8.6630 0.6790 8.9380 1.5430 ;
    LAYER M1 ;
      RECT 1.0390 0.7130 1.1650 0.7630 ;
      RECT 1.0390 0.7630 1.0890 1.0330 ;
      RECT 1.1150 0.5630 1.1650 0.7130 ;
      RECT 1.0230 0.5130 1.1650 0.5630 ;
      RECT 2.9990 0.3880 3.6730 0.4380 ;
      RECT 3.6230 0.4380 3.6730 0.5630 ;
      RECT 3.6230 0.2970 3.6730 0.3880 ;
      RECT 3.4710 0.9670 3.6890 1.0170 ;
      RECT 3.4710 0.3840 3.5210 0.3880 ;
      RECT 3.4710 0.4380 3.5210 0.9670 ;
      RECT 3.4710 1.0170 3.5210 1.1200 ;
      RECT 3.4710 1.1700 3.5210 1.2700 ;
      RECT 2.9990 1.1200 3.5210 1.1700 ;
      RECT 2.3890 0.8580 2.5490 0.9080 ;
      RECT 2.3890 0.9080 2.4390 0.9680 ;
      RECT 1.8590 0.9680 2.4390 1.0180 ;
      RECT 1.3430 0.8540 2.2450 0.9040 ;
      RECT 1.3430 0.9040 1.3930 1.0590 ;
      RECT 1.3430 0.6130 1.3930 0.8540 ;
      RECT 1.3430 1.0590 1.7130 1.1090 ;
      RECT 1.3430 0.5630 1.5450 0.6130 ;
      RECT 1.3430 1.1090 1.3930 1.3370 ;
      RECT 1.4950 0.4070 1.5450 0.5630 ;
      RECT 1.3430 0.4130 1.3930 0.5630 ;
      RECT 4.7630 0.6420 5.2850 0.6920 ;
      RECT 4.1190 0.4500 4.1690 0.7290 ;
      RECT 4.1190 0.7290 4.4850 0.7790 ;
      RECT 4.4350 0.7790 4.4850 1.1790 ;
      RECT 4.7630 0.4500 4.8130 0.6420 ;
      RECT 3.7750 0.4000 4.8130 0.4500 ;
      RECT 3.7760 1.1790 4.4850 1.2290 ;
      RECT 3.7750 0.4500 3.8250 0.5630 ;
      RECT 3.7750 0.2970 3.8250 0.4000 ;
      RECT 3.7760 1.2290 3.8260 1.3530 ;
      RECT 3.6230 0.8670 3.7650 0.9170 ;
      RECT 3.6230 0.6630 3.6730 0.8670 ;
      RECT 3.6230 0.6130 4.0690 0.6630 ;
      RECT 2.7110 0.9200 3.1410 0.9700 ;
      RECT 3.0910 0.8310 3.1410 0.9200 ;
      RECT 2.7110 0.9700 2.7610 1.0340 ;
      RECT 2.7110 0.5050 2.7610 0.9200 ;
      RECT 2.4670 1.4200 3.7730 1.4700 ;
      RECT 1.4790 1.1900 1.8650 1.2400 ;
      RECT 4.0560 1.2790 4.4490 1.3290 ;
      RECT 1.4030 1.3890 1.9410 1.4390 ;
      RECT 3.3230 0.1880 3.9170 0.2380 ;
      RECT 3.3230 0.2380 3.3730 0.2880 ;
      RECT 2.6820 0.2880 3.3730 0.3380 ;
      RECT 2.2950 0.4550 2.3450 0.6130 ;
      RECT 1.8590 0.6130 2.3450 0.6630 ;
      RECT 2.6820 0.3380 2.7320 0.4050 ;
      RECT 2.2950 0.4050 2.7320 0.4550 ;
      RECT 1.1910 0.8130 1.2810 0.8630 ;
      RECT 1.1910 0.8630 1.2410 1.0830 ;
      RECT 1.2310 0.4620 1.2810 0.8130 ;
      RECT 0.4310 1.0830 1.2410 1.1330 ;
      RECT 1.1750 0.4120 1.2810 0.4620 ;
      RECT 1.1910 1.1330 1.2410 1.3540 ;
      RECT 0.4310 0.7980 0.4810 1.0830 ;
      RECT 0.4310 0.7480 0.5210 0.7980 ;
      RECT 0.4310 0.4350 0.5210 0.4850 ;
      RECT 0.4310 0.3720 0.4810 0.4350 ;
      RECT 0.4710 0.4850 0.5210 0.7480 ;
      RECT 5.3370 0.6130 5.8930 0.6630 ;
      RECT 4.5350 0.7920 4.5850 1.3010 ;
      RECT 4.5350 0.5500 4.5850 0.7420 ;
      RECT 4.3070 0.5000 4.5850 0.5500 ;
      RECT 4.3070 0.5500 4.3570 0.6790 ;
      RECT 4.8390 0.7920 4.8890 1.3010 ;
      RECT 5.3370 0.6630 5.3870 0.7420 ;
      RECT 4.5350 0.7420 5.3870 0.7920 ;
      RECT 5.8110 1.1990 7.1090 1.2490 ;
      RECT 3.9340 0.9670 4.0690 1.0170 ;
      RECT 3.9340 0.9160 3.9840 0.9670 ;
      RECT 3.8350 0.8660 3.9840 0.9160 ;
      RECT 2.8470 0.4880 3.4090 0.5380 ;
      RECT 3.3590 0.5380 3.4090 1.0200 ;
      RECT 2.8630 1.0200 3.4090 1.0700 ;
      RECT 2.5990 0.7880 2.6490 1.1200 ;
      RECT 1.5500 0.7380 2.6510 0.7880 ;
      RECT 2.4070 0.5050 2.4570 0.7380 ;
      RECT 2.8630 1.0700 2.9130 1.1200 ;
      RECT 2.0870 1.1200 2.9130 1.1700 ;
      RECT 0.5830 0.6130 1.0290 0.6630 ;
      RECT 0.5830 0.6630 0.6330 1.0040 ;
      RECT 0.5830 0.4130 0.6330 0.6130 ;
      RECT 0.7940 0.0940 1.4910 0.1440 ;
      RECT 4.6110 0.1380 4.6610 0.1700 ;
      RECT 1.7230 0.0880 4.6610 0.1380 ;
      RECT 1.7230 0.1380 1.7730 0.1700 ;
      RECT 6.7990 0.8200 7.3470 0.8700 ;
      RECT 7.1030 0.7090 7.6410 0.7590 ;
      RECT 7.7270 0.6770 7.7770 0.7680 ;
      RECT 7.6870 0.4270 7.7770 0.4620 ;
      RECT 7.7270 0.1260 7.7770 0.4270 ;
      RECT 7.6870 0.6270 7.7770 0.6770 ;
      RECT 7.6870 0.5120 7.7370 0.6270 ;
      RECT 7.4830 0.4770 7.7370 0.5120 ;
      RECT 7.4830 0.4620 7.7770 0.4770 ;
      RECT 7.1030 0.1320 7.3370 0.1820 ;
      RECT 6.3590 1.0620 6.8080 1.1120 ;
      RECT 6.3590 0.6770 6.4090 1.0620 ;
      RECT 6.3190 0.6270 6.4090 0.6770 ;
      RECT 6.3190 0.4770 6.3690 0.6270 ;
      RECT 6.3190 0.4270 6.4090 0.4770 ;
      RECT 6.3590 0.1260 6.4090 0.4270 ;
      RECT 1.0990 1.5240 2.0930 1.5740 ;
      RECT 6.4190 0.5270 7.0170 0.5770 ;
      RECT 6.6630 0.5770 6.7130 0.8840 ;
      RECT 6.6630 0.1260 6.7130 0.5270 ;
      RECT 6.9670 0.5770 7.0170 0.7700 ;
      RECT 6.9670 0.3480 7.0170 0.5270 ;
      RECT 7.3310 1.0620 7.8690 1.1120 ;
      RECT 6.7990 0.2480 7.6410 0.2980 ;
      RECT 3.3770 1.5200 6.8050 1.5700 ;
      RECT 2.6190 1.5200 3.3090 1.5700 ;
      RECT 3.0740 0.6130 3.3090 0.6630 ;
  END
END RDFFSRASX2_LVT

MACRO PMT2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.912 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.8560 0.3590 0.9670 ;
        RECT 0.2790 0.9670 0.3290 1.5550 ;
        RECT 0.2490 0.8310 0.6330 0.8560 ;
        RECT 0.2790 0.8060 0.6330 0.8310 ;
        RECT 0.5830 0.8560 0.6330 1.5550 ;
    END
    ANTENNADIFFAREA 0.1632 ;
    ANTENNAGATEAREA 0.1632 ;
  END S

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 0.9120 1.7020 ;
    END
  END VDD

  PIN D
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 1.4590 0.5110 1.5750 ;
        RECT 0.4310 0.9210 0.4810 1.4590 ;
    END
    ANTENNADIFFAREA 0.0976 ;
  END D

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 0.9120 0.0300 ;
    END
  END VSS

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6590 0.5730 0.7090 ;
        RECT 0.4010 0.5530 0.5110 0.6590 ;
    END
    ANTENNAGATEAREA 0.048 ;
  END G
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.0270 1.7730 ;
    LAYER PO ;
      RECT 0.0610 0.6430 0.0910 1.6050 ;
      RECT 0.2130 0.6430 0.2430 1.6050 ;
      RECT 0.3650 0.6430 0.3950 1.6050 ;
      RECT 0.5170 0.6430 0.5470 1.6050 ;
      RECT 0.6690 0.6430 0.6990 1.6010 ;
      RECT 0.8210 0.6430 0.8510 1.6050 ;
  END
END PMT2_LVT

MACRO PMT3_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.216 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6590 0.8770 0.7090 ;
        RECT 0.4010 0.5530 0.5110 0.6590 ;
    END
    ANTENNAGATEAREA 0.096 ;
  END G

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.2160 0.0300 ;
    END
  END VSS

  PIN D
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 1.5050 0.7850 1.5550 ;
        RECT 0.4010 1.4590 0.5110 1.5050 ;
        RECT 0.4010 1.5550 0.5110 1.5750 ;
        RECT 0.7350 0.9210 0.7850 1.5050 ;
        RECT 0.4310 0.9210 0.4810 1.4590 ;
    END
    ANTENNADIFFAREA 0.1952 ;
  END D

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.2160 1.7020 ;
    END
  END VDD

  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.8680 0.3590 0.9730 ;
        RECT 0.2790 0.9730 0.3290 1.5550 ;
        RECT 0.2490 0.8430 0.9370 0.8680 ;
        RECT 0.2790 0.8180 0.9370 0.8430 ;
        RECT 0.5830 0.8680 0.6330 1.3710 ;
        RECT 0.8870 0.8680 0.9370 1.5550 ;
    END
    ANTENNADIFFAREA 0.2608 ;
    ANTENNAGATEAREA 0.2608 ;
  END S
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.3310 1.7730 ;
    LAYER PO ;
      RECT 0.9730 0.6430 1.0030 1.6050 ;
      RECT 0.5170 0.6430 0.5470 1.6050 ;
      RECT 0.6690 0.6430 0.6990 1.6050 ;
      RECT 0.8210 0.6430 0.8510 1.6050 ;
      RECT 1.1250 0.6430 1.1550 1.6050 ;
      RECT 0.3650 0.6430 0.3950 1.6050 ;
      RECT 0.2130 0.6430 0.2430 1.6050 ;
      RECT 0.0610 0.6430 0.0910 1.6050 ;
  END
END PMT3_LVT

MACRO RDFFARX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.968 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 6.7990 0.9420 8.2660 1.0020 ;
        RECT 8.1560 0.6900 8.2660 0.9420 ;
    END
  END VDDG

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8870 0.3010 6.4410 0.3510 ;
        RECT 6.3310 0.2490 6.4410 0.3010 ;
        RECT 6.3310 0.3510 6.4410 0.3590 ;
        RECT 6.3870 0.3590 6.4370 0.9690 ;
        RECT 5.9030 0.9690 6.4370 1.0190 ;
        RECT 5.9030 1.0190 5.9530 1.3270 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0970 0.9670 1.1810 1.0170 ;
        RECT 0.0970 1.0170 0.2070 1.1190 ;
    END
    ANTENNAGATEAREA 0.018 ;
  END D

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 8.9680 0.0300 ;
        RECT 0.5830 0.0300 0.6330 0.3070 ;
        RECT 7.8790 0.0300 7.9290 0.3120 ;
        RECT 6.8150 0.0300 6.8650 0.2060 ;
        RECT 0.4310 0.0300 0.4810 0.5570 ;
        RECT 5.7510 0.0300 5.8010 0.2410 ;
        RECT 7.5750 0.0300 7.6250 0.2020 ;
        RECT 5.4870 0.0300 5.5370 0.2830 ;
        RECT 0.5830 0.3070 2.3050 0.3570 ;
        RECT 3.1510 0.2830 5.5370 0.3330 ;
        RECT 2.2550 0.3570 2.3050 0.5770 ;
        RECT 1.4950 0.3570 1.5450 0.5580 ;
        RECT 1.7990 0.3570 1.8490 0.5580 ;
        RECT 5.4470 0.3330 5.4970 0.4430 ;
    END
  END VSS

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2480 1.4650 0.4220 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.5990 0.1570 5.6490 0.4010 ;
        RECT 5.5990 0.4010 6.2990 0.4510 ;
        RECT 6.1770 0.4510 6.2990 0.5380 ;
        RECT 6.2490 0.5380 6.2990 0.8590 ;
        RECT 5.5990 0.8590 6.2990 0.9090 ;
        RECT 5.5990 0.9090 5.6490 1.2320 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 8.9680 1.7020 ;
        RECT 0.5430 1.3400 0.5930 1.6420 ;
        RECT 3.8150 1.3400 3.8650 1.6420 ;
        RECT 0.4130 1.2900 5.8010 1.3400 ;
        RECT 3.1670 0.9730 3.2170 1.2900 ;
        RECT 5.7510 0.9590 5.8010 1.2900 ;
    END
  END VDD

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2890 0.8510 3.4440 0.9670 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END RSTB

  PIN RETN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.1210 1.4080 7.5060 1.4580 ;
        RECT 7.3960 1.3130 7.5060 1.4080 ;
    END
    ANTENNAGATEAREA 0.084 ;
  END RETN
  OBS
    LAYER PO ;
      RECT 2.7970 0.0660 2.8270 0.6910 ;
      RECT 2.3410 0.0660 2.3710 0.6370 ;
      RECT 0.9730 0.8390 1.0030 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 4.6210 0.9390 4.6510 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 2.7970 0.8390 2.8270 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6140 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 4.1650 0.9590 4.1950 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 6.1410 0.0670 6.1710 1.6050 ;
      RECT 1.8850 0.9390 1.9150 1.6060 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.7090 0.0660 3.7390 1.6060 ;
      RECT 1.8850 0.0660 1.9150 0.6370 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 0.9730 0.0660 1.0030 0.6910 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 2.3410 0.9390 2.3710 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 4.1650 0.0660 4.1950 0.6910 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 4.6210 0.0660 4.6510 0.7910 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
    LAYER NWELL ;
      RECT -0.1160 1.5430 9.0770 1.7730 ;
      RECT -0.1160 0.6790 6.0340 1.5430 ;
      RECT 8.8020 0.6790 9.0770 1.5430 ;
      RECT 6.4960 0.4910 8.3420 1.0830 ;
    LAYER M1 ;
      RECT 2.7510 0.0920 5.2850 0.1420 ;
      RECT 2.5590 1.0170 2.6090 1.1900 ;
      RECT 2.5190 0.9670 2.6090 1.0170 ;
      RECT 2.5590 1.1900 2.7610 1.2400 ;
      RECT 2.5190 0.8170 2.5690 0.9670 ;
      RECT 2.7110 0.9740 2.7610 1.1900 ;
      RECT 2.5190 0.7670 2.6490 0.8170 ;
      RECT 2.5990 0.5630 2.6490 0.7670 ;
      RECT 2.5590 0.5130 2.7610 0.5630 ;
      RECT 2.5590 0.2770 2.6090 0.5130 ;
      RECT 2.7110 0.2440 2.7610 0.5130 ;
      RECT 2.7110 0.1940 2.8010 0.2440 ;
      RECT 2.7510 0.1420 2.8010 0.1940 ;
      RECT 2.0630 0.8670 2.3450 0.9170 ;
      RECT 2.2950 0.9170 2.3450 1.1270 ;
      RECT 1.1910 1.1270 2.3450 1.1770 ;
      RECT 1.1910 1.1770 1.2410 1.2400 ;
      RECT 1.2410 0.9170 1.2910 1.0660 ;
      RECT 1.1910 0.4130 1.2410 0.8670 ;
      RECT 1.1910 1.0670 1.2910 1.1270 ;
      RECT 1.2310 1.0660 1.2910 1.0670 ;
      RECT 1.1910 0.8670 1.4850 0.9170 ;
      RECT 2.0630 0.6070 2.1130 0.8670 ;
      RECT 2.0630 0.5570 2.1530 0.6070 ;
      RECT 2.1030 0.4130 2.1530 0.5570 ;
      RECT 4.7470 0.7590 6.1970 0.8090 ;
      RECT 5.6750 0.6420 5.7250 0.7590 ;
      RECT 5.2950 0.8090 5.3450 1.2400 ;
      RECT 5.1030 0.5630 5.1530 0.7590 ;
      RECT 5.1030 0.5130 5.3450 0.5630 ;
      RECT 5.2950 0.3830 5.3450 0.5130 ;
      RECT 1.6470 0.9670 2.2450 1.0170 ;
      RECT 1.3430 0.4070 1.3930 0.6190 ;
      RECT 1.6470 1.0170 1.6970 1.0770 ;
      RECT 1.6470 0.6690 1.6970 0.9670 ;
      RECT 1.3430 0.6190 1.6970 0.6690 ;
      RECT 1.6470 0.4070 1.6970 0.6190 ;
      RECT 3.0150 0.5130 3.1050 0.5630 ;
      RECT 3.0550 0.5630 3.1050 0.7670 ;
      RECT 2.9750 0.7670 3.1050 0.8170 ;
      RECT 2.8630 0.2770 3.0650 0.3270 ;
      RECT 2.8630 0.3270 2.9130 0.5560 ;
      RECT 3.0150 0.3270 3.0650 0.5130 ;
      RECT 2.9750 0.8170 3.0250 0.9740 ;
      RECT 2.9750 0.9740 3.0650 1.0240 ;
      RECT 3.0150 1.0240 3.0650 1.1900 ;
      RECT 2.8630 1.1900 3.0650 1.2400 ;
      RECT 2.8630 0.9740 2.9130 1.1900 ;
      RECT 7.7270 0.5890 7.9200 0.6390 ;
      RECT 7.8700 0.5120 7.9200 0.5890 ;
      RECT 7.8700 0.4620 8.0210 0.5120 ;
      RECT 7.8700 0.4120 7.9200 0.4620 ;
      RECT 7.7270 0.3620 7.9200 0.4120 ;
      RECT 7.7270 0.6390 7.7770 0.7820 ;
      RECT 7.7270 0.1260 7.7770 0.3620 ;
      RECT 2.7710 0.6130 3.0050 0.6630 ;
      RECT 0.6430 1.5240 3.0050 1.5740 ;
      RECT 0.7950 0.0940 2.7010 0.1440 ;
      RECT 3.7350 0.7670 3.9770 0.8170 ;
      RECT 3.9270 0.8170 3.9770 1.2400 ;
      RECT 3.7350 0.4530 3.7850 0.7670 ;
      RECT 3.1550 0.4030 3.9770 0.4530 ;
      RECT 3.6230 0.4530 3.6730 0.5770 ;
      RECT 3.9270 0.4530 3.9770 0.5770 ;
      RECT 3.1550 0.4530 3.2050 0.8670 ;
      RECT 3.0750 0.8670 3.2050 0.9170 ;
      RECT 4.0390 0.5130 4.9050 0.5630 ;
      RECT 4.0390 0.5630 4.0890 0.6270 ;
      RECT 3.8350 0.6270 4.0890 0.6770 ;
      RECT 4.0390 0.6770 4.0890 1.0670 ;
      RECT 4.0390 1.0670 4.9050 1.1170 ;
      RECT 4.1390 0.6130 5.0410 0.6630 ;
      RECT 4.9910 0.3830 5.0410 0.6130 ;
      RECT 4.3430 0.6630 4.3930 0.9670 ;
      RECT 4.3430 0.9670 5.0410 1.0170 ;
      RECT 4.9910 1.0170 5.0410 1.2400 ;
      RECT 7.4230 0.4620 7.7170 0.5120 ;
      RECT 7.4230 0.1820 7.4730 0.4620 ;
      RECT 7.4230 0.5120 7.4730 0.6350 ;
      RECT 7.1030 0.1320 7.4730 0.1820 ;
      RECT 7.1030 0.6350 7.4730 0.6850 ;
      RECT 6.9670 0.4940 7.3210 0.5440 ;
      RECT 7.2710 0.3480 7.3210 0.4940 ;
      RECT 6.9670 0.5440 7.0170 0.7820 ;
      RECT 4.2910 1.5280 8.3270 1.5780 ;
      RECT 4.4430 0.7130 4.6770 0.7630 ;
      RECT 8.0310 0.5620 8.3250 0.6120 ;
      RECT 8.1660 0.4120 8.2160 0.5620 ;
      RECT 8.0310 0.3620 8.2160 0.4120 ;
      RECT 8.0310 0.6120 8.0810 0.8320 ;
      RECT 6.8670 0.8320 8.0810 0.8820 ;
      RECT 8.0310 0.1260 8.0810 0.3620 ;
      RECT 6.8670 0.4200 6.9170 0.8320 ;
      RECT 6.8670 0.3700 7.0350 0.4200 ;
      RECT 2.6190 0.8670 2.8730 0.9170 ;
      RECT 0.2790 0.6130 0.7250 0.6630 ;
      RECT 0.6090 0.4630 0.6590 0.6130 ;
      RECT 0.6090 0.4130 1.0130 0.4630 ;
      RECT 0.9630 0.4630 1.0130 0.6800 ;
      RECT 0.2790 0.6630 0.3290 0.9120 ;
      RECT 0.2790 0.4130 0.3290 0.6130 ;
      RECT 0.7190 0.5130 0.8610 0.5630 ;
      RECT 0.8110 0.5630 0.8610 0.7130 ;
      RECT 0.7350 0.7130 0.8610 0.7630 ;
      RECT 0.7350 0.7630 0.7850 0.8670 ;
      RECT 0.7350 0.8670 1.0290 0.9170 ;
      RECT 3.4710 1.0320 3.5640 1.0820 ;
      RECT 3.4710 1.0820 3.5210 1.2400 ;
      RECT 3.5140 0.9170 3.5640 1.0320 ;
      RECT 3.5140 0.8670 3.7650 0.9170 ;
      RECT 3.5140 0.7810 3.5640 0.8670 ;
      RECT 3.4710 0.7310 3.5640 0.7810 ;
      RECT 3.4710 0.5050 3.5210 0.7310 ;
      RECT 1.5490 1.3900 3.7650 1.4400 ;
      RECT 2.1630 0.6670 2.5490 0.7170 ;
      RECT 6.1150 1.2000 7.2610 1.2500 ;
      RECT 5.5750 0.5010 5.8770 0.5510 ;
      RECT 5.8270 0.5510 5.8770 0.6790 ;
      RECT 5.5750 0.5510 5.6250 0.6130 ;
      RECT 5.2030 0.6130 5.6250 0.6630 ;
      RECT 6.6630 1.0620 7.1090 1.1120 ;
      RECT 6.6630 0.1260 6.7130 1.0620 ;
  END
END RDFFARX1_LVT

MACRO RDFFARX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.272 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 7.1030 0.9420 8.5700 1.0020 ;
        RECT 8.4600 0.6900 8.5700 0.9420 ;
    END
  END VDDG

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.7510 0.1490 5.8010 0.4020 ;
        RECT 5.7510 0.4020 6.6030 0.4520 ;
        RECT 6.4810 0.4520 6.6030 0.5120 ;
        RECT 6.5530 0.5120 6.6030 0.8330 ;
        RECT 5.7510 0.8330 6.6030 0.8830 ;
        RECT 5.7510 0.8830 5.8010 1.2240 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0970 0.9670 1.1810 1.0170 ;
        RECT 0.0970 1.0170 0.2070 1.1190 ;
    END
    ANTENNAGATEAREA 0.018 ;
  END D

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.0550 0.2710 6.7530 0.3210 ;
        RECT 6.6330 0.3210 6.7530 0.3600 ;
        RECT 6.6330 0.2500 6.7530 0.2710 ;
        RECT 6.0550 0.1490 6.1050 0.2710 ;
        RECT 6.7030 0.3600 6.7530 0.9330 ;
        RECT 6.6330 0.2470 6.7450 0.2500 ;
        RECT 6.0550 0.9330 6.7530 0.9830 ;
        RECT 6.0550 0.9830 6.1050 1.2240 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 9.2720 0.0300 ;
        RECT 0.5830 0.0300 0.6330 0.3070 ;
        RECT 8.1830 0.0300 8.2330 0.3120 ;
        RECT 5.9030 0.0300 5.9530 0.3200 ;
        RECT 7.1190 0.0300 7.1690 0.2060 ;
        RECT 6.2070 0.0300 6.2570 0.2210 ;
        RECT 0.4310 0.0300 0.4810 0.5570 ;
        RECT 5.5990 0.0300 5.6490 0.4090 ;
        RECT 7.8790 0.0300 7.9290 0.2020 ;
        RECT 5.4870 0.0300 5.5370 0.2830 ;
        RECT 0.5830 0.3070 2.3050 0.3570 ;
        RECT 3.1510 0.2830 5.5370 0.3330 ;
        RECT 2.2550 0.3570 2.3050 0.5770 ;
        RECT 1.4950 0.3570 1.5450 0.5580 ;
        RECT 1.7990 0.3570 1.8490 0.5580 ;
        RECT 5.4470 0.3330 5.4970 0.4430 ;
    END
  END VSS

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 1.4650 0.4220 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 9.2720 1.7020 ;
        RECT 0.5430 1.3400 0.5930 1.6420 ;
        RECT 3.8150 1.3400 3.8650 1.6420 ;
        RECT 0.4130 1.2900 6.2570 1.3400 ;
        RECT 6.2070 1.0530 6.2570 1.2900 ;
        RECT 5.9030 0.9610 5.9530 1.2900 ;
        RECT 5.5990 0.9130 5.6490 1.2900 ;
        RECT 3.1670 0.9730 3.2170 1.2900 ;
    END
  END VDD

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2880 0.8510 3.4440 0.9670 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END RSTB

  PIN RETN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.1210 1.4080 7.8100 1.4580 ;
        RECT 7.6970 1.3130 7.8100 1.4080 ;
    END
    ANTENNAGATEAREA 0.084 ;
  END RETN
  OBS
    LAYER M1 ;
      RECT 6.9670 0.1260 7.0170 1.0620 ;
      RECT 2.7510 0.0920 5.2850 0.1420 ;
      RECT 2.5190 0.7670 2.6490 0.8170 ;
      RECT 2.5990 0.5630 2.6490 0.7670 ;
      RECT 2.5190 0.8170 2.5690 0.9670 ;
      RECT 2.5590 0.5130 2.7610 0.5630 ;
      RECT 2.5190 0.9670 2.6090 1.0170 ;
      RECT 2.5590 0.2770 2.6090 0.5130 ;
      RECT 2.7110 0.2440 2.7610 0.5130 ;
      RECT 2.5590 1.0170 2.6090 1.1900 ;
      RECT 2.7110 0.1940 2.8010 0.2440 ;
      RECT 2.5590 1.1900 2.7610 1.2400 ;
      RECT 2.7510 0.1420 2.8010 0.1940 ;
      RECT 2.7110 0.9740 2.7610 1.1900 ;
      RECT 2.0630 0.8670 2.3450 0.9170 ;
      RECT 2.2950 0.9170 2.3450 1.1270 ;
      RECT 1.1910 1.1270 2.3450 1.1770 ;
      RECT 1.1910 1.1770 1.2410 1.2400 ;
      RECT 1.2410 0.9170 1.2910 1.0660 ;
      RECT 1.1910 0.4130 1.2410 0.8670 ;
      RECT 1.1910 1.0670 1.2910 1.1270 ;
      RECT 1.2310 1.0660 1.2910 1.0670 ;
      RECT 1.1910 0.8670 1.4850 0.9170 ;
      RECT 2.0630 0.6070 2.1130 0.8670 ;
      RECT 2.0630 0.5570 2.1530 0.6070 ;
      RECT 2.1030 0.4130 2.1530 0.5570 ;
      RECT 8.3350 0.5620 8.6290 0.6120 ;
      RECT 8.4700 0.4120 8.5200 0.5620 ;
      RECT 8.3350 0.3620 8.5200 0.4120 ;
      RECT 8.3350 0.6120 8.3850 0.8320 ;
      RECT 7.1710 0.8320 8.3850 0.8820 ;
      RECT 8.3350 0.1260 8.3850 0.3620 ;
      RECT 7.1710 0.4200 7.2210 0.8320 ;
      RECT 7.1710 0.3700 7.3390 0.4200 ;
      RECT 1.6470 0.9670 2.2450 1.0170 ;
      RECT 1.3430 0.4070 1.3930 0.6190 ;
      RECT 1.6470 1.0170 1.6970 1.0770 ;
      RECT 1.6470 0.6690 1.6970 0.9670 ;
      RECT 1.3430 0.6190 1.6970 0.6690 ;
      RECT 1.6470 0.4070 1.6970 0.6190 ;
      RECT 4.7470 0.7130 6.5010 0.7630 ;
      RECT 5.2950 0.7630 5.3450 1.2400 ;
      RECT 5.1030 0.5630 5.1530 0.7130 ;
      RECT 5.1030 0.5130 5.3450 0.5630 ;
      RECT 5.2950 0.3830 5.3450 0.5130 ;
      RECT 5.6750 0.6420 5.7250 0.7130 ;
      RECT 5.8270 0.6420 5.8770 0.7130 ;
      RECT 3.0150 0.5130 3.1050 0.5630 ;
      RECT 3.0550 0.5630 3.1050 0.7670 ;
      RECT 2.9750 0.7670 3.1050 0.8170 ;
      RECT 2.8630 0.2770 3.0650 0.3270 ;
      RECT 2.8630 0.3270 2.9130 0.5560 ;
      RECT 3.0150 0.3270 3.0650 0.5130 ;
      RECT 2.9750 0.8170 3.0250 0.9740 ;
      RECT 2.9750 0.9740 3.0650 1.0240 ;
      RECT 3.0150 1.0240 3.0650 1.1900 ;
      RECT 2.8630 1.1900 3.0650 1.2400 ;
      RECT 2.8630 0.9740 2.9130 1.1900 ;
      RECT 8.0310 0.5890 8.2240 0.6390 ;
      RECT 8.1740 0.5120 8.2240 0.5890 ;
      RECT 8.1740 0.4620 8.3250 0.5120 ;
      RECT 8.1740 0.4120 8.2240 0.4620 ;
      RECT 8.0310 0.3620 8.2240 0.4120 ;
      RECT 8.0310 0.6390 8.0810 0.7430 ;
      RECT 8.0310 0.1260 8.0810 0.3620 ;
      RECT 2.7710 0.6130 3.0050 0.6630 ;
      RECT 0.6430 1.5240 3.0050 1.5740 ;
      RECT 0.7950 0.0940 2.7010 0.1440 ;
      RECT 3.7350 0.7670 3.9770 0.8170 ;
      RECT 3.9270 0.8170 3.9770 1.2400 ;
      RECT 3.7350 0.4530 3.7850 0.7670 ;
      RECT 3.1550 0.4030 3.9770 0.4530 ;
      RECT 3.6230 0.4530 3.6730 0.5770 ;
      RECT 3.9270 0.4530 3.9770 0.5770 ;
      RECT 3.1550 0.4530 3.2050 0.8670 ;
      RECT 3.0750 0.8670 3.2050 0.9170 ;
      RECT 4.0390 0.5130 4.9050 0.5630 ;
      RECT 4.0390 0.5630 4.0890 0.6270 ;
      RECT 3.8350 0.6270 4.0890 0.6770 ;
      RECT 4.0390 0.6770 4.0890 1.0670 ;
      RECT 4.0390 1.0670 4.9050 1.1170 ;
      RECT 4.1390 0.6130 5.0410 0.6630 ;
      RECT 4.9910 0.3830 5.0410 0.6130 ;
      RECT 4.3430 0.6630 4.3930 0.9670 ;
      RECT 4.3430 0.9670 5.0410 1.0170 ;
      RECT 4.9910 1.0170 5.0410 1.2400 ;
      RECT 7.7270 0.4620 8.0210 0.5120 ;
      RECT 7.7270 0.1820 7.7770 0.4620 ;
      RECT 7.7270 0.5120 7.7770 0.6350 ;
      RECT 7.4070 0.1320 7.7770 0.1820 ;
      RECT 7.4070 0.6350 7.7770 0.6850 ;
      RECT 7.2710 0.4940 7.6250 0.5440 ;
      RECT 7.5750 0.3480 7.6250 0.4940 ;
      RECT 7.2710 0.5440 7.3210 0.7720 ;
      RECT 4.2910 1.5280 8.6310 1.5780 ;
      RECT 4.4430 0.7130 4.6770 0.7630 ;
      RECT 2.6190 0.8670 2.8730 0.9170 ;
      RECT 0.2790 0.6130 0.7250 0.6630 ;
      RECT 0.6090 0.4630 0.6590 0.6130 ;
      RECT 0.6090 0.4130 1.0130 0.4630 ;
      RECT 0.9630 0.4630 1.0130 0.6800 ;
      RECT 0.2790 0.6630 0.3290 0.9120 ;
      RECT 0.2790 0.4130 0.3290 0.6130 ;
      RECT 0.7190 0.5130 0.8610 0.5630 ;
      RECT 0.8110 0.5630 0.8610 0.7130 ;
      RECT 0.7350 0.7130 0.8610 0.7630 ;
      RECT 0.7350 0.7630 0.7850 0.8670 ;
      RECT 0.7350 0.8670 1.0290 0.9170 ;
      RECT 3.4710 1.0320 3.5640 1.0820 ;
      RECT 3.4710 1.0820 3.5210 1.2400 ;
      RECT 3.5140 0.9170 3.5640 1.0320 ;
      RECT 3.5140 0.8670 3.7650 0.9170 ;
      RECT 3.5140 0.7810 3.5640 0.8670 ;
      RECT 3.4710 0.7310 3.5640 0.7810 ;
      RECT 3.4710 0.5050 3.5210 0.7310 ;
      RECT 1.5490 1.3900 3.7650 1.4400 ;
      RECT 2.1630 0.6670 2.5490 0.7170 ;
      RECT 6.4190 1.2000 7.5650 1.2500 ;
      RECT 5.5260 0.5200 6.0110 0.5700 ;
      RECT 5.9610 0.5700 6.0110 0.6040 ;
      RECT 5.5260 0.5700 5.5760 0.6130 ;
      RECT 5.9610 0.6040 6.1970 0.6540 ;
      RECT 5.2030 0.6130 5.5760 0.6630 ;
      RECT 6.9670 1.0620 7.4130 1.1120 ;
    LAYER PO ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 2.7970 0.0660 2.8270 0.6910 ;
      RECT 2.3410 0.0660 2.3710 0.6370 ;
      RECT 0.9730 0.8390 1.0030 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 4.6210 0.9390 4.6510 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 2.7970 0.8390 2.8270 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6140 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 4.1650 0.9590 4.1950 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 6.4450 0.0670 6.4750 1.6050 ;
      RECT 1.8850 0.9390 1.9150 1.6060 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.7090 0.0660 3.7390 1.6060 ;
      RECT 1.8850 0.0660 1.9150 0.6370 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 0.9730 0.0660 1.0030 0.6910 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 2.3410 0.9390 2.3710 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 4.1650 0.0660 4.1950 0.6910 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 4.6210 0.0660 4.6510 0.7910 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
    LAYER NWELL ;
      RECT -0.1160 1.5430 9.3810 1.7730 ;
      RECT -0.1160 0.6790 6.3380 1.5430 ;
      RECT 9.1060 0.6790 9.3810 1.5430 ;
      RECT 6.8000 0.4910 8.6460 1.0830 ;
  END
END RDFFARX2_LVT

MACRO RDFFNARX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.968 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 6.7990 0.9420 8.2660 1.0020 ;
        RECT 8.1560 0.6900 8.2660 0.9420 ;
    END
  END VDDG

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.8870 0.3010 6.4410 0.3510 ;
        RECT 6.3280 0.2490 6.4410 0.3010 ;
        RECT 6.3280 0.3510 6.4410 0.3590 ;
        RECT 6.3870 0.3590 6.4370 0.9690 ;
        RECT 5.9030 0.9690 6.4370 1.0190 ;
        RECT 5.9030 1.0190 5.9530 1.3270 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0970 0.9670 1.1810 1.0170 ;
        RECT 0.0970 1.0170 0.2070 1.1190 ;
    END
    ANTENNAGATEAREA 0.018 ;
  END D

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 8.9680 0.0300 ;
        RECT 7.8790 0.0300 7.9290 0.3120 ;
        RECT 6.8150 0.0300 6.8650 0.2060 ;
        RECT 5.7510 0.0300 5.8010 0.2410 ;
        RECT 7.5750 0.0300 7.6250 0.2020 ;
        RECT 5.4870 0.0300 5.5370 0.2830 ;
        RECT 0.3910 0.0300 0.4410 0.3060 ;
        RECT 3.1510 0.2830 5.5370 0.3330 ;
        RECT 0.3910 0.3060 0.4810 0.3070 ;
        RECT 5.4470 0.3330 5.4970 0.4430 ;
        RECT 0.3910 0.3070 2.3050 0.3570 ;
        RECT 0.4310 0.3570 0.4810 0.5570 ;
        RECT 2.2550 0.3570 2.3050 0.5770 ;
        RECT 1.4950 0.3570 1.5450 0.5580 ;
        RECT 1.7990 0.3570 1.8490 0.5580 ;
    END
  END VSS

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2480 1.4650 0.4220 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.5990 0.1570 5.6490 0.4010 ;
        RECT 5.5990 0.4010 6.2990 0.4510 ;
        RECT 6.1770 0.4510 6.2990 0.5380 ;
        RECT 6.2490 0.5380 6.2990 0.8590 ;
        RECT 5.5990 0.8590 6.2990 0.9090 ;
        RECT 5.5990 0.9090 5.6490 1.2320 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 8.9680 1.7020 ;
        RECT 0.5430 1.3400 0.5930 1.6420 ;
        RECT 3.8150 1.3400 3.8650 1.6420 ;
        RECT 0.4130 1.2900 5.8010 1.3400 ;
        RECT 3.1670 0.9730 3.2170 1.2900 ;
        RECT 5.7510 0.9590 5.8010 1.2900 ;
    END
  END VDD

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2880 0.8510 3.4440 0.9670 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END RSTB

  PIN RETN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.1210 1.4080 7.5060 1.4580 ;
        RECT 7.3910 1.3130 7.5060 1.4080 ;
    END
    ANTENNAGATEAREA 0.084 ;
  END RETN
  OBS
    LAYER PO ;
      RECT 4.6210 0.9390 4.6510 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 2.7970 0.8390 2.8270 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6140 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 4.1650 0.9590 4.1950 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 6.1410 0.0670 6.1710 1.6050 ;
      RECT 1.8850 0.9390 1.9150 1.6060 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.7090 0.0660 3.7390 1.6060 ;
      RECT 1.8850 0.0660 1.9150 0.6370 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 0.9730 0.0660 1.0030 0.6910 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 2.3410 0.9390 2.3710 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 4.1650 0.0660 4.1950 0.6910 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 4.6210 0.0660 4.6510 0.7910 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 2.7970 0.0660 2.8270 0.6910 ;
      RECT 2.3410 0.0660 2.3710 0.6370 ;
      RECT 0.9730 0.8390 1.0030 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
    LAYER NWELL ;
      RECT -0.1160 1.5430 9.0770 1.7730 ;
      RECT -0.1160 0.6790 6.0340 1.5430 ;
      RECT 8.8020 0.6790 9.0770 1.5430 ;
      RECT 6.4960 0.4910 8.3420 1.0830 ;
    LAYER M1 ;
      RECT 2.7510 0.0920 5.2850 0.1420 ;
      RECT 2.7110 0.9740 2.7610 1.1900 ;
      RECT 2.5590 1.1900 2.7610 1.2400 ;
      RECT 2.5590 1.0170 2.6090 1.1900 ;
      RECT 2.5190 0.9670 2.6090 1.0170 ;
      RECT 2.5190 0.8170 2.5690 0.9670 ;
      RECT 2.5190 0.7670 2.6490 0.8170 ;
      RECT 2.5990 0.5630 2.6490 0.7670 ;
      RECT 2.5590 0.5130 2.7610 0.5630 ;
      RECT 2.5590 0.2770 2.6090 0.5130 ;
      RECT 2.7110 0.2440 2.7610 0.5130 ;
      RECT 2.7110 0.1940 2.8010 0.2440 ;
      RECT 2.7510 0.1420 2.8010 0.1940 ;
      RECT 3.0150 0.5130 3.1050 0.5630 ;
      RECT 3.0550 0.5630 3.1050 0.7670 ;
      RECT 2.9750 0.7670 3.1050 0.8170 ;
      RECT 2.8630 0.2770 3.0650 0.3270 ;
      RECT 2.8630 0.3270 2.9130 0.5560 ;
      RECT 3.0150 0.3270 3.0650 0.5130 ;
      RECT 2.9750 0.8170 3.0250 0.9740 ;
      RECT 2.9750 0.9740 3.0650 1.0240 ;
      RECT 3.0150 1.0240 3.0650 1.1900 ;
      RECT 2.8630 1.1900 3.0650 1.2400 ;
      RECT 2.8630 0.9740 2.9130 1.1900 ;
      RECT 1.6470 0.9670 2.2450 1.0170 ;
      RECT 1.3430 0.4070 1.3930 0.6190 ;
      RECT 1.6470 1.0170 1.6970 1.0770 ;
      RECT 1.6470 0.6690 1.6970 0.9670 ;
      RECT 1.3430 0.6190 1.6970 0.6690 ;
      RECT 1.6470 0.4070 1.6970 0.6190 ;
      RECT 7.7270 0.5890 7.9200 0.6390 ;
      RECT 7.8700 0.5120 7.9200 0.5890 ;
      RECT 7.8700 0.4620 8.0210 0.5120 ;
      RECT 7.8700 0.4120 7.9200 0.4620 ;
      RECT 7.7270 0.3620 7.9200 0.4120 ;
      RECT 7.7270 0.6390 7.7770 0.7750 ;
      RECT 7.7270 0.1260 7.7770 0.3620 ;
      RECT 2.7710 0.6130 3.0050 0.6630 ;
      RECT 2.0630 0.8670 2.3450 0.9170 ;
      RECT 2.2950 0.9170 2.3450 1.1270 ;
      RECT 1.1910 1.1270 2.3450 1.1770 ;
      RECT 1.1910 1.1770 1.2410 1.2400 ;
      RECT 1.2410 0.9170 1.2910 1.0660 ;
      RECT 1.1910 0.4130 1.2410 0.8670 ;
      RECT 1.1910 1.0670 1.2910 1.1270 ;
      RECT 1.2310 1.0660 1.2910 1.0670 ;
      RECT 1.1910 0.8670 1.4850 0.9170 ;
      RECT 2.0630 0.6070 2.1130 0.8670 ;
      RECT 2.0630 0.5570 2.1530 0.6070 ;
      RECT 2.1030 0.4130 2.1530 0.5570 ;
      RECT 0.7950 1.5240 3.0050 1.5740 ;
      RECT 0.4910 0.0940 2.7010 0.1440 ;
      RECT 3.7350 0.7670 3.9770 0.8170 ;
      RECT 3.9270 0.8170 3.9770 1.2400 ;
      RECT 3.7350 0.4530 3.7850 0.7670 ;
      RECT 3.1550 0.4030 3.9770 0.4530 ;
      RECT 3.6230 0.4530 3.6730 0.5770 ;
      RECT 3.9270 0.4530 3.9770 0.5770 ;
      RECT 3.1550 0.4530 3.2050 0.8670 ;
      RECT 3.0750 0.8670 3.2050 0.9170 ;
      RECT 4.0390 0.5130 4.9050 0.5630 ;
      RECT 4.0390 0.5630 4.0890 0.6270 ;
      RECT 3.8350 0.6270 4.0890 0.6770 ;
      RECT 4.0390 0.6770 4.0890 1.0670 ;
      RECT 4.0390 1.0670 4.9050 1.1170 ;
      RECT 4.1390 0.6130 5.0410 0.6630 ;
      RECT 4.9910 0.3830 5.0410 0.6130 ;
      RECT 4.3430 0.6630 4.3930 0.9670 ;
      RECT 4.3430 0.9670 5.0410 1.0170 ;
      RECT 4.9910 1.0170 5.0410 1.2400 ;
      RECT 7.4230 0.4620 7.7170 0.5120 ;
      RECT 7.4230 0.1820 7.4730 0.4620 ;
      RECT 7.4230 0.5120 7.4730 0.6350 ;
      RECT 7.1030 0.1320 7.4730 0.1820 ;
      RECT 7.1030 0.6350 7.4730 0.6850 ;
      RECT 6.9670 0.4940 7.3210 0.5440 ;
      RECT 7.2710 0.3480 7.3210 0.4940 ;
      RECT 6.9670 0.5440 7.0170 0.7520 ;
      RECT 4.7470 0.7590 6.1970 0.8090 ;
      RECT 5.6750 0.6420 5.7250 0.7590 ;
      RECT 5.2950 0.8090 5.3450 1.2400 ;
      RECT 5.1030 0.5630 5.1530 0.7590 ;
      RECT 5.1030 0.5130 5.3450 0.5630 ;
      RECT 5.2950 0.3830 5.3450 0.5130 ;
      RECT 4.2910 1.5280 8.3270 1.5780 ;
      RECT 4.4430 0.7130 4.6770 0.7630 ;
      RECT 8.0310 0.5620 8.3250 0.6120 ;
      RECT 8.1660 0.4120 8.2160 0.5620 ;
      RECT 8.0310 0.3620 8.2160 0.4120 ;
      RECT 8.0310 0.6120 8.0810 0.8320 ;
      RECT 6.8670 0.8320 8.0810 0.8820 ;
      RECT 8.0310 0.1260 8.0810 0.3620 ;
      RECT 6.8670 0.4200 6.9170 0.8320 ;
      RECT 6.8670 0.3700 7.0350 0.4200 ;
      RECT 2.6190 0.8670 2.8730 0.9170 ;
      RECT 0.2790 0.6130 0.7250 0.6630 ;
      RECT 0.2790 0.8670 1.0290 0.9170 ;
      RECT 0.2790 0.4130 0.3290 0.6130 ;
      RECT 0.2790 0.6630 0.3290 0.8670 ;
      RECT 0.7190 0.5130 0.8610 0.5630 ;
      RECT 0.8110 0.5630 0.8610 0.6130 ;
      RECT 0.8110 0.6130 1.0300 0.6630 ;
      RECT 0.8110 0.6630 0.8610 0.7540 ;
      RECT 0.7170 0.7540 0.8610 0.8040 ;
      RECT 3.4710 1.0320 3.5640 1.0820 ;
      RECT 3.4710 1.0820 3.5210 1.2400 ;
      RECT 3.5140 0.9170 3.5640 1.0320 ;
      RECT 3.5140 0.8670 3.7650 0.9170 ;
      RECT 3.5140 0.7810 3.5640 0.8670 ;
      RECT 3.4710 0.7310 3.5640 0.7810 ;
      RECT 3.4710 0.5050 3.5210 0.7310 ;
      RECT 1.5490 1.3900 3.7650 1.4400 ;
      RECT 2.1630 0.6670 2.5490 0.7170 ;
      RECT 6.1150 1.2000 7.2610 1.2500 ;
      RECT 5.5750 0.5010 5.8770 0.5510 ;
      RECT 5.8270 0.5510 5.8770 0.6790 ;
      RECT 5.5750 0.5510 5.6250 0.6130 ;
      RECT 5.2030 0.6130 5.6250 0.6630 ;
      RECT 6.6630 1.0620 7.1090 1.1120 ;
      RECT 6.6630 0.1260 6.7130 1.0620 ;
  END
END RDFFNARX1_LVT

MACRO RDFFNARX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.272 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 7.1030 0.9420 8.5700 1.0020 ;
        RECT 8.4600 0.6900 8.5700 0.9420 ;
    END
  END VDDG

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.4810 0.3990 6.5930 0.4020 ;
        RECT 5.7510 0.4020 6.6030 0.4520 ;
        RECT 5.7510 0.1490 5.8010 0.4020 ;
        RECT 6.4810 0.4520 6.6030 0.5120 ;
        RECT 6.5530 0.5120 6.6030 0.8330 ;
        RECT 5.7510 0.8330 6.6030 0.8830 ;
        RECT 5.7510 0.8830 5.8010 1.2240 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0970 0.9670 1.1810 1.0170 ;
        RECT 0.0970 1.0170 0.2070 1.1190 ;
    END
    ANTENNAGATEAREA 0.018 ;
  END D

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 9.2720 0.0300 ;
        RECT 8.1830 0.0300 8.2330 0.3120 ;
        RECT 7.1190 0.0300 7.1690 0.2060 ;
        RECT 5.9030 0.0300 5.9530 0.3200 ;
        RECT 6.2070 0.0300 6.2570 0.2210 ;
        RECT 5.5990 0.0300 5.6490 0.4090 ;
        RECT 7.8790 0.0300 7.9290 0.2020 ;
        RECT 5.4870 0.0300 5.5370 0.2830 ;
        RECT 0.3910 0.0300 0.4410 0.3060 ;
        RECT 3.1510 0.2830 5.5370 0.3330 ;
        RECT 0.3910 0.3060 0.4810 0.3070 ;
        RECT 5.4470 0.3330 5.4970 0.4430 ;
        RECT 0.3910 0.3070 2.3050 0.3570 ;
        RECT 0.4310 0.3570 0.4810 0.5570 ;
        RECT 2.2550 0.3570 2.3050 0.5770 ;
        RECT 1.4950 0.3570 1.5450 0.5580 ;
        RECT 1.7990 0.3570 1.8490 0.5580 ;
    END
  END VSS

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2470 1.4650 0.4220 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.0550 0.1490 6.1050 0.2710 ;
        RECT 6.0550 0.2710 6.7530 0.3210 ;
        RECT 6.6330 0.2450 6.7530 0.2710 ;
        RECT 6.6330 0.3210 6.7530 0.3600 ;
        RECT 6.7030 0.3600 6.7530 0.9330 ;
        RECT 6.0550 0.9330 6.7530 0.9830 ;
        RECT 6.0550 0.9830 6.1050 1.2240 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 9.2720 1.7020 ;
        RECT 0.5430 1.3400 0.5930 1.6420 ;
        RECT 3.8150 1.3400 3.8650 1.6420 ;
        RECT 0.4130 1.2900 6.2570 1.3400 ;
        RECT 6.2070 1.0530 6.2570 1.2900 ;
        RECT 5.9030 0.9610 5.9530 1.2900 ;
        RECT 5.5990 0.9130 5.6490 1.2900 ;
        RECT 3.1670 0.9730 3.2170 1.2900 ;
    END
  END VDD

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2880 0.8510 3.4440 0.9670 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END RSTB

  PIN RETN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.1210 1.4080 7.8100 1.4580 ;
        RECT 7.6930 1.3130 7.8100 1.4080 ;
    END
    ANTENNAGATEAREA 0.084 ;
  END RETN
  OBS
    LAYER PO ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 2.7970 0.0660 2.8270 0.6910 ;
      RECT 2.3410 0.0660 2.3710 0.6370 ;
      RECT 0.9730 0.8390 1.0030 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 4.6210 0.9390 4.6510 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 2.7970 0.8390 2.8270 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6140 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 4.1650 0.9590 4.1950 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 6.4450 0.0670 6.4750 1.6050 ;
      RECT 1.8850 0.9390 1.9150 1.6060 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.7090 0.0660 3.7390 1.6060 ;
      RECT 1.8850 0.0660 1.9150 0.6370 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 0.9730 0.0660 1.0030 0.6910 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 9.1810 0.0660 9.2110 1.6060 ;
      RECT 2.3410 0.9390 2.3710 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 9.0290 0.0660 9.0590 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 4.1650 0.0660 4.1950 0.6910 ;
      RECT 8.8770 0.0660 8.9070 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 8.5730 0.0660 8.6030 1.6060 ;
      RECT 4.6210 0.0660 4.6510 0.7910 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 8.7250 0.0660 8.7550 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
    LAYER NWELL ;
      RECT -0.1160 1.5430 9.3810 1.7730 ;
      RECT -0.1160 0.6790 6.3380 1.5430 ;
      RECT 9.1060 0.6790 9.3810 1.5430 ;
      RECT 6.8000 0.4910 8.6460 1.0830 ;
    LAYER M1 ;
      RECT 5.9610 0.6040 6.1970 0.6540 ;
      RECT 5.9610 0.5700 6.0110 0.6040 ;
      RECT 5.5260 0.5200 6.0110 0.5700 ;
      RECT 5.5260 0.5700 5.5760 0.6130 ;
      RECT 5.2030 0.6130 5.5760 0.6630 ;
      RECT 6.9670 1.0620 7.4130 1.1120 ;
      RECT 6.9670 0.1260 7.0170 1.0620 ;
      RECT 2.7510 0.0920 5.2850 0.1420 ;
      RECT 2.7510 0.1420 2.8010 0.1940 ;
      RECT 2.7110 0.1940 2.8010 0.2440 ;
      RECT 2.7110 0.2440 2.7610 0.5130 ;
      RECT 2.5590 0.5130 2.7610 0.5630 ;
      RECT 2.5590 0.2770 2.6090 0.5130 ;
      RECT 2.5990 0.5630 2.6490 0.7670 ;
      RECT 2.5190 0.7670 2.6490 0.8170 ;
      RECT 2.5190 0.8170 2.5690 0.9670 ;
      RECT 2.5190 0.9670 2.6090 1.0170 ;
      RECT 2.5590 1.0170 2.6090 1.1900 ;
      RECT 2.5590 1.1900 2.7610 1.2400 ;
      RECT 2.7110 0.9740 2.7610 1.1900 ;
      RECT 2.0630 0.8670 2.3450 0.9170 ;
      RECT 2.2950 0.9170 2.3450 1.1270 ;
      RECT 1.1910 1.1270 2.3450 1.1770 ;
      RECT 1.1910 1.1770 1.2410 1.2400 ;
      RECT 1.2410 0.9170 1.2910 1.0660 ;
      RECT 1.1910 0.4130 1.2410 0.8670 ;
      RECT 1.1910 1.0670 1.2910 1.1270 ;
      RECT 1.2310 1.0660 1.2910 1.0670 ;
      RECT 1.1910 0.8670 1.4850 0.9170 ;
      RECT 2.0630 0.6070 2.1130 0.8670 ;
      RECT 2.0630 0.5570 2.1530 0.6070 ;
      RECT 2.1030 0.4130 2.1530 0.5570 ;
      RECT 8.3350 0.5620 8.6290 0.6120 ;
      RECT 8.4700 0.4120 8.5200 0.5620 ;
      RECT 8.3350 0.3620 8.5200 0.4120 ;
      RECT 8.3350 0.6120 8.3850 0.8320 ;
      RECT 7.1710 0.8320 8.3850 0.8820 ;
      RECT 8.3350 0.1260 8.3850 0.3620 ;
      RECT 7.1710 0.4200 7.2210 0.8320 ;
      RECT 7.1710 0.3700 7.3390 0.4200 ;
      RECT 1.6470 0.9670 2.2450 1.0170 ;
      RECT 1.3430 0.4070 1.3930 0.6190 ;
      RECT 1.6470 1.0170 1.6970 1.0770 ;
      RECT 1.6470 0.6690 1.6970 0.9670 ;
      RECT 1.3430 0.6190 1.6970 0.6690 ;
      RECT 1.6470 0.4070 1.6970 0.6190 ;
      RECT 3.0150 0.5130 3.1050 0.5630 ;
      RECT 3.0550 0.5630 3.1050 0.7670 ;
      RECT 2.9750 0.7670 3.1050 0.8170 ;
      RECT 2.8630 0.2770 3.0650 0.3270 ;
      RECT 2.8630 0.3270 2.9130 0.5560 ;
      RECT 3.0150 0.3270 3.0650 0.5130 ;
      RECT 2.9750 0.8170 3.0250 0.9740 ;
      RECT 2.9750 0.9740 3.0650 1.0240 ;
      RECT 3.0150 1.0240 3.0650 1.1900 ;
      RECT 2.8630 1.1900 3.0650 1.2400 ;
      RECT 2.8630 0.9740 2.9130 1.1900 ;
      RECT 8.0310 0.5890 8.2240 0.6390 ;
      RECT 8.1740 0.5120 8.2240 0.5890 ;
      RECT 8.1740 0.4620 8.3250 0.5120 ;
      RECT 8.1740 0.4120 8.2240 0.4620 ;
      RECT 8.0310 0.3620 8.2240 0.4120 ;
      RECT 8.0310 0.6390 8.0810 0.7280 ;
      RECT 8.0310 0.1260 8.0810 0.3620 ;
      RECT 2.7710 0.6130 3.0050 0.6630 ;
      RECT 0.7950 1.5240 3.0050 1.5740 ;
      RECT 0.4910 0.0940 2.7010 0.1440 ;
      RECT 3.7350 0.7670 3.9770 0.8170 ;
      RECT 3.9270 0.8170 3.9770 1.2400 ;
      RECT 3.7350 0.4530 3.7850 0.7670 ;
      RECT 3.1550 0.4030 3.9770 0.4530 ;
      RECT 3.6230 0.4530 3.6730 0.5770 ;
      RECT 3.9270 0.4530 3.9770 0.5770 ;
      RECT 3.1550 0.4530 3.2050 0.8670 ;
      RECT 3.0750 0.8670 3.2050 0.9170 ;
      RECT 4.0390 0.5130 4.9050 0.5630 ;
      RECT 4.0390 0.5630 4.0890 0.6270 ;
      RECT 3.8350 0.6270 4.0890 0.6770 ;
      RECT 4.0390 0.6770 4.0890 1.0670 ;
      RECT 4.0390 1.0670 4.9050 1.1170 ;
      RECT 4.1390 0.6130 5.0410 0.6630 ;
      RECT 4.9910 0.3830 5.0410 0.6130 ;
      RECT 4.3430 0.6630 4.3930 0.9670 ;
      RECT 4.3430 0.9670 5.0410 1.0170 ;
      RECT 4.9910 1.0170 5.0410 1.2400 ;
      RECT 7.7270 0.4620 8.0210 0.5120 ;
      RECT 7.7270 0.1820 7.7770 0.4620 ;
      RECT 7.7270 0.5120 7.7770 0.6350 ;
      RECT 7.4070 0.1320 7.7770 0.1820 ;
      RECT 7.4070 0.6350 7.7770 0.6850 ;
      RECT 7.2710 0.4940 7.6250 0.5440 ;
      RECT 7.5750 0.3480 7.6250 0.4940 ;
      RECT 7.2710 0.5440 7.3210 0.7730 ;
      RECT 4.2910 1.5280 8.6310 1.5780 ;
      RECT 4.4430 0.7130 4.6770 0.7630 ;
      RECT 2.6190 0.8670 2.8730 0.9170 ;
      RECT 0.2790 0.6130 0.7250 0.6630 ;
      RECT 0.2790 0.8670 1.0290 0.9170 ;
      RECT 0.2790 0.4130 0.3290 0.6130 ;
      RECT 0.2790 0.6630 0.3290 0.8670 ;
      RECT 0.7190 0.5130 0.8610 0.5630 ;
      RECT 0.8110 0.5630 0.8610 0.6130 ;
      RECT 0.8110 0.6130 1.0300 0.6630 ;
      RECT 0.8110 0.6630 0.8610 0.7540 ;
      RECT 0.7170 0.7540 0.8610 0.8040 ;
      RECT 3.4710 1.0320 3.5640 1.0820 ;
      RECT 3.4710 1.0820 3.5210 1.2400 ;
      RECT 3.5140 0.9170 3.5640 1.0320 ;
      RECT 3.5140 0.8670 3.7650 0.9170 ;
      RECT 3.5140 0.7810 3.5640 0.8670 ;
      RECT 3.4710 0.7310 3.5640 0.7810 ;
      RECT 3.4710 0.5050 3.5210 0.7310 ;
      RECT 1.5490 1.3900 3.7650 1.4400 ;
      RECT 2.1630 0.6670 2.5490 0.7170 ;
      RECT 6.4190 1.2000 7.5650 1.2500 ;
      RECT 4.7470 0.7130 6.5010 0.7630 ;
      RECT 5.2950 0.7630 5.3450 1.2400 ;
      RECT 5.1030 0.5630 5.1530 0.7130 ;
      RECT 5.1030 0.5130 5.3450 0.5630 ;
      RECT 5.2950 0.3830 5.3450 0.5130 ;
      RECT 5.6750 0.6420 5.7250 0.7130 ;
      RECT 5.8270 0.6420 5.8770 0.7130 ;
  END
END RDFFNARX2_LVT

MACRO RDFFNSRARX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.208 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.4650 0.7250 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.4210 0.6630 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 8.2080 1.7020 ;
        RECT 0.2790 1.1310 0.3290 1.6420 ;
        RECT 2.1430 1.2700 2.1930 1.6420 ;
        RECT 6.2470 1.4540 6.2970 1.6420 ;
        RECT 0.4480 1.2940 0.4980 1.6420 ;
        RECT 1.9340 1.2200 3.0810 1.2700 ;
        RECT 3.7750 1.4040 6.2970 1.4540 ;
        RECT 0.4480 1.2440 0.9530 1.2940 ;
        RECT 3.7750 1.2790 3.8250 1.4040 ;
        RECT 4.8390 0.9590 4.8890 1.4040 ;
        RECT 4.3830 0.9530 4.4330 1.4040 ;
    END
  END VDD

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6870 0.4010 5.3870 0.4510 ;
        RECT 4.6870 0.1570 4.7370 0.4010 ;
        RECT 5.2650 0.4510 5.3870 0.5380 ;
        RECT 5.3370 0.5380 5.3870 0.8590 ;
        RECT 4.6870 0.8590 5.3870 0.9090 ;
        RECT 4.6870 0.9090 4.7370 1.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.9910 0.9690 5.5250 1.0190 ;
        RECT 5.4750 0.3510 5.5250 0.9690 ;
        RECT 4.9910 1.0190 5.2230 1.1290 ;
        RECT 4.9750 0.3010 5.5250 0.3510 ;
        RECT 4.9910 1.1290 5.0410 1.3270 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 8.2080 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.2720 ;
        RECT 4.8390 0.0300 4.8890 0.2410 ;
        RECT 6.8150 0.0300 6.8650 0.1980 ;
        RECT 7.2710 0.0300 7.3210 0.4260 ;
        RECT 5.9030 0.0300 5.9530 0.4260 ;
        RECT 4.5590 0.0300 4.6090 0.3000 ;
        RECT 0.2790 0.2720 2.1530 0.3220 ;
        RECT 3.7590 0.3000 4.6090 0.3500 ;
        RECT 1.9510 0.3220 2.0010 0.5570 ;
        RECT 0.7350 0.3220 0.7850 0.5570 ;
        RECT 0.8870 0.3220 0.9370 0.5570 ;
        RECT 2.1030 0.3220 2.1530 0.3470 ;
        RECT 0.2790 0.3220 0.3290 0.4050 ;
        RECT 2.1030 0.2380 2.1530 0.2720 ;
        RECT 2.1030 0.1880 3.0810 0.2380 ;
        RECT 2.4070 0.2380 2.4570 0.3490 ;
    END
  END VSS

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6150 0.0970 3.8650 0.1380 ;
        RECT 1.6150 0.1380 1.7730 0.2100 ;
        RECT 3.8150 0.1380 3.8650 0.2000 ;
        RECT 1.7230 0.0880 3.8650 0.0970 ;
        RECT 3.8150 0.2000 4.3570 0.2500 ;
        RECT 4.3070 0.0880 4.3570 0.2000 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.3900 0.2490 7.5050 0.3590 ;
        RECT 7.4040 0.3590 7.4540 0.5270 ;
        RECT 7.1790 0.5270 7.4540 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6810 0.7040 2.8370 0.7310 ;
        RECT 2.6810 0.7310 3.1410 0.7810 ;
        RECT 2.7870 0.5970 2.8370 0.7040 ;
        RECT 2.6810 0.7810 2.8370 0.8150 ;
        RECT 3.0910 0.7810 3.1410 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 5.8870 0.9420 7.5050 1.0020 ;
        RECT 7.3950 0.6900 7.5050 0.9420 ;
        RECT 7.2710 0.6270 7.3210 0.9420 ;
    END
  END VDDG
  OBS
    LAYER PO ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 2.7970 0.0660 2.8270 0.6910 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 1.8850 0.9390 1.9150 1.6060 ;
      RECT 5.2290 0.0670 5.2590 1.6050 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 3.1010 0.8390 3.1310 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 3.8610 0.0660 3.8910 0.6910 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 3.7090 0.0660 3.7390 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 1.2770 0.8400 1.3070 1.6060 ;
      RECT 3.8610 0.9390 3.8910 1.6060 ;
      RECT 3.5570 0.0660 3.5870 0.6370 ;
      RECT 1.2770 0.0660 1.3070 0.6370 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 1.8850 0.0660 1.9150 0.6910 ;
      RECT 3.1010 0.0660 3.1310 0.6910 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 2.7970 0.8920 2.8270 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
      RECT 3.5570 0.8390 3.5870 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
    LAYER NWELL ;
      RECT 5.5840 0.4910 7.5950 1.0830 ;
      RECT -0.1150 1.5430 8.3300 1.7730 ;
      RECT -0.1150 0.6790 5.1220 1.5430 ;
      RECT 8.0550 0.6790 8.3300 1.5430 ;
    LAYER M1 ;
      RECT 3.3190 0.9670 3.5370 1.0170 ;
      RECT 3.3190 0.4380 3.3690 0.9670 ;
      RECT 3.3190 1.0170 3.3690 1.1200 ;
      RECT 2.8470 0.3880 3.5210 0.4380 ;
      RECT 3.4710 0.4380 3.5210 0.5630 ;
      RECT 3.4710 0.2970 3.5210 0.3880 ;
      RECT 3.3190 0.3840 3.3690 0.3880 ;
      RECT 3.3190 1.1700 3.3690 1.2700 ;
      RECT 2.8470 1.1200 3.3690 1.1700 ;
      RECT 2.2970 0.8580 2.3970 0.9080 ;
      RECT 2.2970 0.9080 2.3470 0.9680 ;
      RECT 1.8590 0.9680 2.3470 1.0180 ;
      RECT 1.3430 0.8540 2.2450 0.9040 ;
      RECT 1.3430 0.9040 1.3930 1.0590 ;
      RECT 1.3430 0.6130 1.3930 0.8540 ;
      RECT 1.3430 1.0590 1.7130 1.1090 ;
      RECT 1.3430 0.5630 1.5450 0.6130 ;
      RECT 1.3430 1.1090 1.3930 1.3370 ;
      RECT 1.4950 0.4070 1.5450 0.5630 ;
      RECT 1.3430 0.4130 1.3930 0.5630 ;
      RECT 4.4590 0.6420 4.8130 0.6920 ;
      RECT 4.7630 0.5970 4.8130 0.6420 ;
      RECT 3.9940 0.4500 4.0440 0.7290 ;
      RECT 3.9940 0.7290 4.1810 0.7790 ;
      RECT 4.1310 0.7790 4.1810 1.1790 ;
      RECT 3.6240 1.1790 4.1810 1.2290 ;
      RECT 4.4590 0.4500 4.5090 0.6420 ;
      RECT 3.6230 0.4000 4.5090 0.4500 ;
      RECT 3.6230 0.4500 3.6730 0.5630 ;
      RECT 3.6230 0.2970 3.6730 0.4000 ;
      RECT 3.6240 1.2290 3.6740 1.3530 ;
      RECT 3.1710 0.1880 3.7650 0.2380 ;
      RECT 3.1710 0.2380 3.2210 0.2880 ;
      RECT 2.5300 0.2880 3.2210 0.3380 ;
      RECT 2.1230 0.4550 2.1730 0.6130 ;
      RECT 1.8590 0.6130 2.1730 0.6630 ;
      RECT 2.5300 0.3380 2.5800 0.4050 ;
      RECT 2.1230 0.4050 2.5800 0.4550 ;
      RECT 4.8630 0.6130 5.2850 0.6630 ;
      RECT 4.2310 0.8090 4.2810 1.3010 ;
      RECT 4.2310 0.6780 4.2810 0.7590 ;
      RECT 4.1390 0.6280 4.2810 0.6780 ;
      RECT 4.2310 0.5000 4.2810 0.6280 ;
      RECT 4.5350 0.8090 4.5850 1.3010 ;
      RECT 4.8630 0.6630 4.9130 0.7590 ;
      RECT 4.2310 0.7590 4.9130 0.8090 ;
      RECT 5.2030 1.1990 6.5010 1.2490 ;
      RECT 3.4710 0.8670 3.6130 0.9170 ;
      RECT 3.4710 0.6630 3.5210 0.8670 ;
      RECT 3.4710 0.6130 3.9170 0.6630 ;
      RECT 3.7820 0.9670 3.9170 1.0170 ;
      RECT 3.7820 0.9160 3.8320 0.9670 ;
      RECT 3.6830 0.8660 3.8320 0.9160 ;
      RECT 3.2070 0.5380 3.2570 1.0200 ;
      RECT 2.6950 0.5070 3.2570 0.5380 ;
      RECT 2.7110 1.0200 3.2570 1.0700 ;
      RECT 2.6950 0.4880 3.2560 0.5070 ;
      RECT 2.4470 0.7880 2.4970 1.1200 ;
      RECT 1.5500 0.7380 2.4990 0.7880 ;
      RECT 2.2550 0.5050 2.3050 0.7380 ;
      RECT 2.7110 1.0700 2.7610 1.1200 ;
      RECT 2.2340 1.1200 2.7610 1.1700 ;
      RECT 1.1910 0.8130 1.2810 0.8630 ;
      RECT 1.2310 0.4620 1.2810 0.8130 ;
      RECT 1.1910 0.8630 1.2410 1.0830 ;
      RECT 1.1750 0.4120 1.2810 0.4620 ;
      RECT 0.4310 1.0830 1.2410 1.1330 ;
      RECT 1.1910 1.1330 1.2410 1.3540 ;
      RECT 0.4310 0.7980 0.4810 1.0830 ;
      RECT 0.4310 0.7480 0.5210 0.7980 ;
      RECT 0.4310 0.4350 0.5210 0.4850 ;
      RECT 0.4310 0.3720 0.4810 0.4350 ;
      RECT 0.4710 0.4850 0.5210 0.7480 ;
      RECT 0.5830 0.6130 1.0290 0.6630 ;
      RECT 0.5830 0.6630 0.6330 1.0040 ;
      RECT 0.5830 0.4130 0.6330 0.6130 ;
      RECT 6.1910 0.8200 6.7390 0.8700 ;
      RECT 6.4950 0.7090 7.0330 0.7590 ;
      RECT 7.1190 0.6770 7.1690 0.7680 ;
      RECT 7.0790 0.4270 7.1690 0.4620 ;
      RECT 7.1190 0.1260 7.1690 0.4270 ;
      RECT 7.0790 0.6270 7.1690 0.6770 ;
      RECT 7.0790 0.5120 7.1290 0.6270 ;
      RECT 6.8750 0.4770 7.1290 0.5120 ;
      RECT 6.8750 0.4620 7.1690 0.4770 ;
      RECT 6.4950 0.1320 6.7290 0.1820 ;
      RECT 5.7510 1.0620 6.2000 1.1120 ;
      RECT 5.7510 0.6770 5.8010 1.0620 ;
      RECT 5.7110 0.6270 5.8010 0.6770 ;
      RECT 5.7110 0.4770 5.7610 0.6270 ;
      RECT 5.7110 0.4270 5.8010 0.4770 ;
      RECT 5.7510 0.1260 5.8010 0.4270 ;
      RECT 5.8110 0.5270 6.4090 0.5770 ;
      RECT 6.0550 0.5770 6.1050 0.8540 ;
      RECT 6.0550 0.1260 6.1050 0.5270 ;
      RECT 6.3590 0.5770 6.4090 0.7700 ;
      RECT 6.3590 0.3480 6.4090 0.5270 ;
      RECT 3.9870 0.0940 4.2210 0.1440 ;
      RECT 6.7230 1.0700 7.2610 1.1200 ;
      RECT 6.1910 0.2480 7.0330 0.2980 ;
      RECT 3.2250 1.5200 6.1970 1.5700 ;
      RECT 0.7950 1.5240 2.0930 1.5740 ;
      RECT 2.4670 1.5200 3.1570 1.5700 ;
      RECT 2.9220 0.6130 3.1570 0.6630 ;
      RECT 2.5590 0.9200 2.9890 0.9700 ;
      RECT 2.9390 0.8310 2.9890 0.9200 ;
      RECT 2.5590 0.9700 2.6090 1.0340 ;
      RECT 2.5590 0.5050 2.6090 0.9200 ;
      RECT 2.3150 1.4200 3.6210 1.4700 ;
      RECT 1.4790 1.1900 1.8650 1.2400 ;
      RECT 1.4030 1.3890 1.9410 1.4390 ;
      RECT 1.0980 0.0940 1.4910 0.1440 ;
      RECT 1.0390 0.7130 1.1650 0.7630 ;
      RECT 1.0390 0.7630 1.0890 1.0330 ;
      RECT 1.1150 0.5630 1.1650 0.7130 ;
      RECT 1.0230 0.5130 1.1650 0.5630 ;
  END
END RDFFNSRARX1_LVT

MACRO RDFFNSRARX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.512 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 6.1910 0.9420 7.8090 1.0020 ;
        RECT 7.6990 0.6900 7.8090 0.9420 ;
        RECT 7.5750 0.6270 7.6250 0.9420 ;
    END
  END VDDG

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6810 0.7030 2.8370 0.7310 ;
        RECT 2.6810 0.7310 3.1410 0.7810 ;
        RECT 2.7870 0.5970 2.8370 0.7030 ;
        RECT 2.6810 0.7810 2.8370 0.8150 ;
        RECT 3.0910 0.7810 3.1410 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.6950 0.2490 7.8090 0.3590 ;
        RECT 7.7080 0.3590 7.7580 0.5270 ;
        RECT 7.4830 0.5270 7.7580 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6150 0.1410 1.7730 0.2100 ;
        RECT 1.6150 0.0970 3.8650 0.1410 ;
        RECT 3.8150 0.1410 3.8650 0.2000 ;
        RECT 1.7230 0.0910 3.8650 0.0970 ;
        RECT 3.8150 0.2000 4.3570 0.2500 ;
        RECT 4.3070 0.0880 4.3570 0.2000 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 8.5120 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.2720 ;
        RECT 7.5750 0.0300 7.6250 0.4260 ;
        RECT 5.2950 0.0300 5.3450 0.2200 ;
        RECT 4.6870 0.0300 4.7370 0.4080 ;
        RECT 6.2070 0.0300 6.2570 0.4260 ;
        RECT 7.1190 0.0300 7.1690 0.1980 ;
        RECT 4.9910 0.0300 5.0410 0.3190 ;
        RECT 4.5590 0.0300 4.6090 0.3000 ;
        RECT 0.2790 0.2720 2.1530 0.3220 ;
        RECT 3.7590 0.3000 4.6090 0.3500 ;
        RECT 0.7350 0.3220 0.7850 0.5570 ;
        RECT 1.9510 0.3220 2.0010 0.5570 ;
        RECT 0.8870 0.3220 0.9370 0.5570 ;
        RECT 2.1030 0.3220 2.1530 0.3470 ;
        RECT 0.2790 0.3220 0.3290 0.4050 ;
        RECT 2.1030 0.2470 2.1530 0.2720 ;
        RECT 2.1030 0.1970 3.0810 0.2470 ;
        RECT 2.4070 0.2470 2.4570 0.3490 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 8.5120 1.7020 ;
        RECT 0.2790 1.1310 0.3290 1.6420 ;
        RECT 6.5510 1.4540 6.6010 1.6420 ;
        RECT 2.1430 1.2700 2.1930 1.6420 ;
        RECT 0.4480 1.2940 0.4980 1.6420 ;
        RECT 3.7750 1.4040 6.6010 1.4540 ;
        RECT 1.9340 1.2200 3.0810 1.2700 ;
        RECT 0.4480 1.2440 0.9530 1.2940 ;
        RECT 3.7750 1.2790 3.8250 1.4040 ;
        RECT 4.6870 0.9120 4.7370 1.4040 ;
        RECT 5.2950 1.0520 5.3450 1.4040 ;
        RECT 4.9910 0.9600 5.0410 1.4040 ;
        RECT 4.3830 0.9530 4.4330 1.4040 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.4210 0.6630 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.4650 0.7250 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.8390 0.1480 4.8890 0.4010 ;
        RECT 4.8390 0.4010 5.6910 0.4510 ;
        RECT 5.5690 0.4510 5.6910 0.5110 ;
        RECT 5.6410 0.5110 5.6910 0.8320 ;
        RECT 4.8390 0.8320 5.6910 0.8820 ;
        RECT 4.8390 0.8820 4.8890 1.3180 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.1430 0.2700 5.8410 0.3200 ;
        RECT 5.7200 0.3200 5.8410 0.3590 ;
        RECT 5.7200 0.2490 5.8410 0.2700 ;
        RECT 5.1430 0.1480 5.1930 0.2700 ;
        RECT 5.7910 0.3590 5.8410 0.9320 ;
        RECT 5.1430 0.9320 5.8410 0.9820 ;
        RECT 5.1430 0.9820 5.1930 1.3260 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q
  OBS
    LAYER PO ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 1.2770 0.0660 1.3070 0.6370 ;
      RECT 3.5570 0.0660 3.5870 0.6370 ;
      RECT 1.2770 0.8400 1.3070 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 3.8610 0.0660 3.8910 0.6910 ;
      RECT 5.5330 0.0670 5.5630 1.6050 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 5.3810 0.0680 5.4110 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 3.7090 0.0660 3.7390 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 2.7970 0.8920 2.8270 1.6060 ;
      RECT 3.5570 0.8390 3.5870 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 1.8850 0.0660 1.9150 0.6910 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 2.7970 0.0660 2.8270 0.6910 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 1.8850 0.9390 1.9150 1.6060 ;
      RECT 3.1010 0.0660 3.1310 0.6910 ;
      RECT 3.8610 0.9390 3.8910 1.6060 ;
      RECT 3.1010 0.8390 3.1310 1.6060 ;
    LAYER NWELL ;
      RECT -0.1150 0.6790 5.4260 1.5430 ;
      RECT -0.1150 1.5430 8.6290 1.7730 ;
      RECT 8.3590 0.6790 8.6290 1.5430 ;
      RECT 5.8880 0.4910 7.8990 1.0830 ;
    LAYER M1 ;
      RECT 1.0390 0.7130 1.1650 0.7630 ;
      RECT 1.0390 0.7630 1.0890 1.0330 ;
      RECT 1.1150 0.5630 1.1650 0.7130 ;
      RECT 1.0230 0.5130 1.1650 0.5630 ;
      RECT 2.8470 0.3970 3.5210 0.4470 ;
      RECT 3.4710 0.4470 3.5210 0.5630 ;
      RECT 3.4710 0.2970 3.5210 0.3970 ;
      RECT 3.3190 0.3840 3.3690 0.3970 ;
      RECT 3.3190 0.4470 3.3690 0.9670 ;
      RECT 3.3190 0.9670 3.5370 1.0170 ;
      RECT 3.3190 1.0170 3.3690 1.1200 ;
      RECT 3.3190 1.1700 3.3690 1.2700 ;
      RECT 2.8470 1.1200 3.3690 1.1700 ;
      RECT 1.8590 0.9680 2.3470 1.0180 ;
      RECT 2.2970 0.9080 2.3470 0.9680 ;
      RECT 2.2970 0.8580 2.3970 0.9080 ;
      RECT 1.3430 0.8540 2.2450 0.9040 ;
      RECT 1.3430 0.6130 1.3930 0.8540 ;
      RECT 1.3430 0.9040 1.3930 1.0590 ;
      RECT 1.3430 0.5630 1.5450 0.6130 ;
      RECT 1.3430 1.0590 1.7130 1.1090 ;
      RECT 1.3430 0.4130 1.3930 0.5630 ;
      RECT 1.4950 0.4070 1.5450 0.5630 ;
      RECT 1.3430 1.1090 1.3930 1.3370 ;
      RECT 4.4410 0.6320 4.9810 0.6820 ;
      RECT 3.6230 0.4500 3.6730 0.5630 ;
      RECT 3.6230 0.2970 3.6730 0.4000 ;
      RECT 3.6240 1.2290 3.6740 1.3530 ;
      RECT 3.9940 0.4500 4.0440 0.7290 ;
      RECT 3.9940 0.7290 4.1810 0.7790 ;
      RECT 4.1310 0.7790 4.1810 1.1790 ;
      RECT 3.6240 1.1790 4.1810 1.2290 ;
      RECT 4.4590 0.4500 4.5090 0.6320 ;
      RECT 3.6230 0.4000 4.5090 0.4500 ;
      RECT 2.9220 0.6130 3.1570 0.6630 ;
      RECT 3.1710 0.1910 3.7650 0.2410 ;
      RECT 2.1230 0.4550 2.1730 0.6130 ;
      RECT 1.8590 0.6130 2.1730 0.6630 ;
      RECT 3.1710 0.2410 3.2210 0.2970 ;
      RECT 2.5300 0.3470 2.5800 0.4050 ;
      RECT 2.1230 0.4050 2.5800 0.4550 ;
      RECT 2.5300 0.2970 3.2210 0.3470 ;
      RECT 3.4710 0.6130 3.9170 0.6630 ;
      RECT 3.4710 0.6630 3.5210 0.8670 ;
      RECT 3.4710 0.8670 3.6130 0.9170 ;
      RECT 1.1910 0.8130 1.2810 0.8630 ;
      RECT 1.2310 0.4620 1.2810 0.8130 ;
      RECT 1.1910 0.8630 1.2410 1.0830 ;
      RECT 1.1750 0.4120 1.2810 0.4620 ;
      RECT 0.4310 1.0830 1.2410 1.1330 ;
      RECT 1.1910 1.1330 1.2410 1.3540 ;
      RECT 0.4310 0.7980 0.4810 1.0830 ;
      RECT 0.4310 0.7480 0.5210 0.7980 ;
      RECT 0.4310 0.4350 0.5210 0.4850 ;
      RECT 0.4310 0.3720 0.4810 0.4350 ;
      RECT 0.4710 0.4850 0.5210 0.7480 ;
      RECT 0.5830 0.6130 1.0290 0.6630 ;
      RECT 0.5830 0.6630 0.6330 1.0040 ;
      RECT 0.5830 0.4130 0.6330 0.6130 ;
      RECT 2.5590 0.9200 2.9890 0.9700 ;
      RECT 2.9390 0.8310 2.9890 0.9200 ;
      RECT 2.5590 0.9700 2.6090 1.0340 ;
      RECT 2.5590 0.5050 2.6090 0.9200 ;
      RECT 3.2070 0.5470 3.2570 1.0200 ;
      RECT 2.7110 1.0200 3.2570 1.0700 ;
      RECT 2.6950 0.4970 3.2560 0.5070 ;
      RECT 2.6950 0.5070 3.2570 0.5470 ;
      RECT 2.4470 0.7880 2.4970 1.1200 ;
      RECT 1.5500 0.7380 2.4990 0.7880 ;
      RECT 2.2550 0.5050 2.3050 0.7380 ;
      RECT 2.7110 1.0700 2.7610 1.1200 ;
      RECT 2.2340 1.1200 2.7610 1.1700 ;
      RECT 5.0470 0.6130 5.5890 0.6630 ;
      RECT 5.0470 0.6630 5.0970 0.7320 ;
      RECT 4.2310 0.7320 5.0970 0.7820 ;
      RECT 4.2310 0.7820 4.2810 1.3010 ;
      RECT 4.2310 0.6780 4.2810 0.7320 ;
      RECT 4.1390 0.6280 4.2810 0.6780 ;
      RECT 4.2310 0.5000 4.2810 0.6280 ;
      RECT 4.5350 0.7820 4.5850 1.3010 ;
      RECT 6.0550 1.0790 6.5040 1.1290 ;
      RECT 6.0550 0.6770 6.1050 1.0790 ;
      RECT 6.0150 0.6270 6.1050 0.6770 ;
      RECT 6.0150 0.4770 6.0650 0.6270 ;
      RECT 6.0150 0.4270 6.1050 0.4770 ;
      RECT 6.0550 0.1260 6.1050 0.4270 ;
      RECT 7.4230 0.6770 7.4730 0.7680 ;
      RECT 7.3830 0.4270 7.4730 0.4620 ;
      RECT 7.4230 0.1260 7.4730 0.4270 ;
      RECT 7.3830 0.6270 7.4730 0.6770 ;
      RECT 7.3830 0.5120 7.4330 0.6270 ;
      RECT 7.1790 0.4770 7.4330 0.5120 ;
      RECT 7.1790 0.4620 7.4730 0.4770 ;
      RECT 5.5070 1.1990 6.8050 1.2490 ;
      RECT 0.7950 1.5240 2.0930 1.5740 ;
      RECT 2.3150 1.4200 3.6210 1.4700 ;
      RECT 3.2250 1.5200 6.5010 1.5700 ;
      RECT 1.0980 0.0940 1.4910 0.1440 ;
      RECT 6.1150 0.5270 6.7130 0.5770 ;
      RECT 6.6630 0.5770 6.7130 0.7700 ;
      RECT 6.6630 0.3480 6.7130 0.5270 ;
      RECT 6.3590 0.5770 6.4090 0.8850 ;
      RECT 6.3590 0.1260 6.4090 0.5270 ;
      RECT 6.7990 0.7090 7.3370 0.7590 ;
      RECT 6.4950 0.8200 7.0430 0.8700 ;
      RECT 6.4950 0.2480 7.3370 0.2980 ;
      RECT 3.9870 0.0940 4.2210 0.1440 ;
      RECT 2.4670 1.5200 3.1570 1.5700 ;
      RECT 7.0270 1.0780 7.5650 1.1280 ;
      RECT 1.4030 1.3890 1.9410 1.4390 ;
      RECT 1.4790 1.1900 1.8650 1.2400 ;
      RECT 3.6830 0.8660 3.8320 0.9160 ;
      RECT 3.7820 0.9160 3.8320 0.9670 ;
      RECT 3.7820 0.9670 3.9170 1.0170 ;
      RECT 6.7990 0.1320 7.0330 0.1820 ;
  END
END RDFFNSRARX2_LVT

MACRO RDFFNSRASRNX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.36 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.4210 0.6630 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 8.3600 1.7020 ;
        RECT 0.2790 1.1310 0.3290 1.6420 ;
        RECT 2.1430 1.2700 2.1930 1.6420 ;
        RECT 0.4310 1.2940 0.4810 1.6420 ;
        RECT 6.3990 1.4540 6.4490 1.6420 ;
        RECT 1.9340 1.2200 3.2330 1.2700 ;
        RECT 0.4310 1.2440 0.9530 1.2940 ;
        RECT 3.9270 1.4040 6.4490 1.4540 ;
        RECT 3.9270 1.2790 3.9770 1.4040 ;
        RECT 5.1430 1.0520 5.1930 1.4040 ;
        RECT 4.6870 0.9530 4.7370 1.4040 ;
    END
  END VDD

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.9910 0.4010 5.5390 0.4510 ;
        RECT 4.9910 0.1570 5.0410 0.4010 ;
        RECT 5.4170 0.4510 5.5390 0.5380 ;
        RECT 5.4890 0.5380 5.5390 0.9520 ;
        RECT 4.9910 0.9520 5.5390 1.0020 ;
        RECT 4.9910 0.9510 5.0410 0.9520 ;
        RECT 4.9910 1.0020 5.0410 1.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 8.3600 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.2720 ;
        RECT 5.1430 0.0300 5.1930 0.2410 ;
        RECT 6.9670 0.0300 7.0170 0.1980 ;
        RECT 7.4230 0.0300 7.4730 0.4260 ;
        RECT 6.0550 0.0300 6.1050 0.4260 ;
        RECT 4.8630 0.0300 4.9130 0.3220 ;
        RECT 0.2790 0.2720 2.1530 0.3220 ;
        RECT 3.9110 0.3220 4.9130 0.3720 ;
        RECT 1.9510 0.3220 2.0010 0.5570 ;
        RECT 0.7350 0.3220 0.7850 0.5570 ;
        RECT 0.8870 0.3220 0.9370 0.5570 ;
        RECT 2.1030 0.3220 2.1530 0.5330 ;
        RECT 0.2790 0.3220 0.3290 0.4050 ;
        RECT 2.1030 0.2470 2.1530 0.2720 ;
        RECT 2.1030 0.1970 3.2330 0.2470 ;
        RECT 2.5590 0.2470 2.6090 0.3490 ;
    END
  END VSS

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.1550 0.8570 4.3110 0.9750 ;
        RECT 4.1550 0.9750 4.2050 1.0790 ;
        RECT 3.6230 1.0790 4.2050 1.1290 ;
        RECT 3.6230 1.1290 3.6730 1.3200 ;
        RECT 2.3310 1.3200 3.6730 1.3700 ;
        RECT 2.3310 1.3700 2.3810 1.4550 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7230 0.0900 4.6610 0.0960 ;
        RECT 1.6150 0.0960 4.6610 0.1400 ;
        RECT 1.6150 0.1400 1.7730 0.2220 ;
        RECT 4.6110 0.1400 4.6610 0.1720 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.4650 0.7250 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.5440 0.2490 7.6570 0.3590 ;
        RECT 7.5560 0.3590 7.6060 0.4980 ;
        RECT 7.3310 0.4980 7.6060 0.5480 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8330 0.7020 2.9890 0.7310 ;
        RECT 2.8330 0.7310 3.2930 0.7810 ;
        RECT 2.9390 0.5970 2.9890 0.7020 ;
        RECT 2.8330 0.7810 2.9890 0.8150 ;
        RECT 3.2430 0.7810 3.2930 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 6.0390 0.9420 7.6570 1.0020 ;
        RECT 7.5470 0.6900 7.6570 0.9420 ;
        RECT 7.4230 0.6270 7.4730 0.9420 ;
    END
  END VDDG
  OBS
    LAYER PO ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 2.9490 0.0660 2.9790 0.6910 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 1.8850 0.9390 1.9150 1.6060 ;
      RECT 5.3810 0.0670 5.4110 1.6050 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 3.2530 0.8390 3.2830 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 4.0130 0.0660 4.0430 0.7540 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 1.2770 0.8400 1.3070 1.6060 ;
      RECT 4.0130 0.9390 4.0430 1.6060 ;
      RECT 3.7090 0.0660 3.7390 0.6370 ;
      RECT 1.2770 0.0660 1.3070 0.6370 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 1.8850 0.0660 1.9150 0.6910 ;
      RECT 3.2530 0.0660 3.2830 0.6910 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 2.9490 0.8920 2.9790 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 3.7090 0.8390 3.7390 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
    LAYER NWELL ;
      RECT 5.7360 0.4910 7.7470 1.0830 ;
      RECT -0.1150 1.5430 8.4820 1.7730 ;
      RECT -0.1150 0.6790 5.2740 1.5430 ;
      RECT 8.2070 0.6790 8.4820 1.5430 ;
    LAYER M1 ;
      RECT 2.9990 0.3970 3.6730 0.4470 ;
      RECT 3.6230 0.4470 3.6730 0.5630 ;
      RECT 3.6230 0.2970 3.6730 0.3970 ;
      RECT 3.4710 0.9670 3.6890 1.0170 ;
      RECT 3.4710 0.4470 3.5210 0.9670 ;
      RECT 3.4710 1.0170 3.5210 1.1200 ;
      RECT 3.4710 1.1700 3.5210 1.2700 ;
      RECT 2.9990 1.1200 3.5210 1.1700 ;
      RECT 2.3890 0.8580 2.5490 0.9080 ;
      RECT 2.3890 0.9080 2.4390 0.9680 ;
      RECT 1.8590 0.9680 2.4390 1.0180 ;
      RECT 1.3430 0.8540 2.2450 0.9040 ;
      RECT 1.3430 0.9040 1.3930 1.0590 ;
      RECT 1.3430 0.6130 1.3930 0.8540 ;
      RECT 1.3430 1.0590 1.7130 1.1090 ;
      RECT 1.3430 0.5630 1.5450 0.6130 ;
      RECT 1.3430 1.1090 1.3930 1.3370 ;
      RECT 1.4950 0.4070 1.5450 0.5630 ;
      RECT 1.3430 0.4130 1.3930 0.5630 ;
      RECT 4.7630 0.6770 5.1170 0.7270 ;
      RECT 5.0670 0.6420 5.1170 0.6770 ;
      RECT 4.1190 0.4920 4.1690 0.7570 ;
      RECT 4.4350 0.8070 4.4850 1.1790 ;
      RECT 4.7630 0.4920 4.8130 0.6770 ;
      RECT 3.7750 0.4420 4.8130 0.4920 ;
      RECT 3.7760 1.1790 4.4850 1.2290 ;
      RECT 4.1190 0.7570 4.4850 0.8070 ;
      RECT 3.7750 0.4920 3.8250 0.5630 ;
      RECT 3.7750 0.2970 3.8250 0.4420 ;
      RECT 3.7760 1.2290 3.8260 1.3530 ;
      RECT 0.7950 1.5240 2.0930 1.5740 ;
      RECT 1.1910 0.8130 1.2810 0.8630 ;
      RECT 1.1910 0.8630 1.2410 1.0830 ;
      RECT 1.2310 0.4620 1.2810 0.8130 ;
      RECT 0.4310 1.0830 1.2410 1.1330 ;
      RECT 1.1750 0.4120 1.2810 0.4620 ;
      RECT 1.1910 1.1330 1.2410 1.3540 ;
      RECT 0.4310 0.7980 0.4810 1.0830 ;
      RECT 0.4310 0.7480 0.5210 0.7980 ;
      RECT 0.4310 0.4350 0.5210 0.4850 ;
      RECT 0.4310 0.3720 0.4810 0.4350 ;
      RECT 0.4710 0.4850 0.5210 0.7480 ;
      RECT 3.3230 0.1910 3.9170 0.2410 ;
      RECT 3.3230 0.2410 3.3730 0.2970 ;
      RECT 2.6820 0.2970 3.3730 0.3470 ;
      RECT 2.2950 0.4550 2.3450 0.6130 ;
      RECT 1.8590 0.6130 2.3450 0.6630 ;
      RECT 2.6820 0.3470 2.7320 0.4050 ;
      RECT 2.2950 0.4050 2.7320 0.4550 ;
      RECT 5.1670 0.6130 5.4370 0.6630 ;
      RECT 4.5350 0.9010 4.5850 1.3010 ;
      RECT 4.5350 0.6070 4.5850 0.8510 ;
      RECT 4.3070 0.5570 4.5850 0.6070 ;
      RECT 4.3070 0.6070 4.3570 0.7070 ;
      RECT 4.5350 0.5420 4.5850 0.5570 ;
      RECT 4.8390 0.9010 4.8890 1.3010 ;
      RECT 5.1670 0.6630 5.2170 0.8510 ;
      RECT 4.5350 0.8510 5.2170 0.9010 ;
      RECT 5.3550 1.1990 6.6530 1.2490 ;
      RECT 3.6230 0.8670 3.7650 0.9170 ;
      RECT 3.6230 0.7220 3.6730 0.8670 ;
      RECT 3.6230 0.6720 4.0690 0.7220 ;
      RECT 3.9340 0.9670 4.0690 1.0170 ;
      RECT 3.9340 0.9160 3.9840 0.9670 ;
      RECT 3.8350 0.8660 3.9840 0.9160 ;
      RECT 2.8470 0.4970 3.4080 0.5070 ;
      RECT 3.3590 0.5470 3.4090 1.0200 ;
      RECT 2.8630 1.0200 3.4090 1.0700 ;
      RECT 2.8470 0.5070 3.4090 0.5470 ;
      RECT 2.5990 0.7880 2.6490 1.1200 ;
      RECT 1.5500 0.7380 2.6510 0.7880 ;
      RECT 2.4070 0.5050 2.4570 0.7380 ;
      RECT 2.8630 1.0700 2.9130 1.1200 ;
      RECT 2.0870 1.1200 2.9130 1.1700 ;
      RECT 0.5830 0.6130 1.0290 0.6630 ;
      RECT 0.5830 0.6630 0.6330 1.0040 ;
      RECT 0.5830 0.4130 0.6330 0.6130 ;
      RECT 6.3430 0.8200 6.8910 0.8700 ;
      RECT 6.6470 0.7090 7.1850 0.7590 ;
      RECT 7.2310 0.6270 7.3210 0.6770 ;
      RECT 7.2710 0.6770 7.3210 0.7680 ;
      RECT 7.2310 0.3870 7.3210 0.4370 ;
      RECT 7.2710 0.1260 7.3210 0.3870 ;
      RECT 7.2310 0.5120 7.2810 0.6270 ;
      RECT 7.0270 0.4620 7.2810 0.5120 ;
      RECT 7.2310 0.4370 7.2810 0.4620 ;
      RECT 6.6470 0.1320 6.8810 0.1820 ;
      RECT 5.9030 1.0690 6.3520 1.1190 ;
      RECT 5.9030 0.6770 5.9530 1.0690 ;
      RECT 5.8630 0.6270 5.9530 0.6770 ;
      RECT 5.8630 0.4770 5.9130 0.6270 ;
      RECT 5.8630 0.4270 5.9530 0.4770 ;
      RECT 5.9030 0.1260 5.9530 0.4270 ;
      RECT 5.9630 0.5270 6.5610 0.5770 ;
      RECT 6.2070 0.5770 6.2570 0.8790 ;
      RECT 6.2070 0.1260 6.2570 0.5270 ;
      RECT 6.5110 0.5770 6.5610 0.7700 ;
      RECT 6.5110 0.3480 6.5610 0.5270 ;
      RECT 6.8750 1.0650 7.4130 1.1150 ;
      RECT 6.3430 0.2480 7.1850 0.2980 ;
      RECT 3.3770 1.5200 6.3490 1.5700 ;
      RECT 1.0980 0.0940 1.4910 0.1440 ;
      RECT 2.6190 1.5200 3.3090 1.5700 ;
      RECT 3.0740 0.6130 3.3090 0.6630 ;
      RECT 2.7110 0.9200 3.1410 0.9700 ;
      RECT 3.0910 0.8310 3.1410 0.9200 ;
      RECT 2.7110 0.9700 2.7610 1.0340 ;
      RECT 2.7110 0.5050 2.7610 0.9200 ;
      RECT 2.4670 1.4200 3.7730 1.4700 ;
      RECT 1.4790 1.1900 1.8650 1.2400 ;
      RECT 4.0560 1.2870 4.4490 1.3370 ;
      RECT 1.4030 1.3890 1.9410 1.4390 ;
      RECT 1.0390 0.7130 1.1650 0.7630 ;
      RECT 1.0390 0.7630 1.0890 1.0330 ;
      RECT 1.1150 0.5630 1.1650 0.7130 ;
      RECT 1.0230 0.5130 1.1650 0.5630 ;
  END
END RDFFNSRASRNX1_LVT

MACRO RDFFNSRASRNX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.512 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.4210 0.6630 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 8.5120 1.7020 ;
        RECT 0.2790 1.1310 0.3290 1.6420 ;
        RECT 2.1430 1.2700 2.1930 1.6420 ;
        RECT 0.4310 1.2940 0.4810 1.6420 ;
        RECT 6.5510 1.4540 6.6010 1.6420 ;
        RECT 1.9340 1.2200 3.2330 1.2700 ;
        RECT 0.4310 1.2440 0.9530 1.2940 ;
        RECT 3.9270 1.4040 6.6010 1.4540 ;
        RECT 3.9270 1.2790 3.9770 1.4040 ;
        RECT 5.1430 0.9590 5.1930 1.4040 ;
        RECT 4.6870 0.9530 4.7370 1.4040 ;
    END
  END VDD

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.9910 0.4010 5.6910 0.4510 ;
        RECT 4.9910 0.1570 5.0410 0.4010 ;
        RECT 5.5690 0.4510 5.6910 0.5110 ;
        RECT 5.2950 0.1570 5.3450 0.4010 ;
        RECT 5.6410 0.5110 5.6910 0.8590 ;
        RECT 4.9910 0.8590 5.6910 0.9090 ;
        RECT 4.9910 0.9090 5.0410 1.3090 ;
        RECT 5.2950 0.9090 5.3450 1.3090 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END QN

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 8.5120 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.2670 ;
        RECT 5.1430 0.0300 5.1930 0.2410 ;
        RECT 7.1190 0.0300 7.1690 0.1980 ;
        RECT 7.5750 0.0300 7.6250 0.4260 ;
        RECT 6.2070 0.0300 6.2570 0.4260 ;
        RECT 4.8630 0.0300 4.9130 0.2880 ;
        RECT 0.2790 0.2670 2.1530 0.3170 ;
        RECT 3.9110 0.2880 4.9130 0.3380 ;
        RECT 1.9510 0.3170 2.0010 0.5570 ;
        RECT 0.7350 0.3170 0.7850 0.5570 ;
        RECT 0.8870 0.3170 0.9370 0.5570 ;
        RECT 2.1030 0.3170 2.1530 0.5330 ;
        RECT 0.2790 0.3170 0.3290 0.4050 ;
        RECT 2.1030 0.2380 2.1530 0.2670 ;
        RECT 2.1030 0.1880 3.2330 0.2380 ;
        RECT 2.5590 0.2380 2.6090 0.3490 ;
    END
  END VSS

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.1550 0.8570 4.3110 0.9750 ;
        RECT 4.1550 0.9750 4.2050 1.0790 ;
        RECT 3.6230 1.0790 4.2050 1.1290 ;
        RECT 3.6230 1.1290 3.6730 1.3200 ;
        RECT 2.3310 1.3200 3.6730 1.3700 ;
        RECT 2.3310 1.3700 2.3810 1.4550 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6150 0.0880 4.6610 0.1380 ;
        RECT 1.6150 0.1380 1.7730 0.2100 ;
        RECT 4.6110 0.1380 4.6610 0.1700 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.4650 0.7250 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.6940 0.2490 7.8090 0.3590 ;
        RECT 7.7080 0.3590 7.7580 0.5270 ;
        RECT 7.4830 0.5270 7.7580 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8330 0.7050 2.9890 0.7310 ;
        RECT 2.8330 0.7310 3.2930 0.7810 ;
        RECT 2.9390 0.5970 2.9890 0.7050 ;
        RECT 2.8330 0.7810 2.9890 0.8150 ;
        RECT 3.2430 0.7810 3.2930 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 6.1910 0.9420 7.8090 1.0020 ;
        RECT 7.6990 0.6900 7.8090 0.9420 ;
        RECT 7.5750 0.6270 7.6250 0.9420 ;
    END
  END VDDG
  OBS
    LAYER PO ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 2.9490 0.0660 2.9790 0.6910 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 1.8850 0.9390 1.9150 1.6060 ;
      RECT 5.5330 0.0670 5.5630 1.6050 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 3.2530 0.8390 3.2830 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 4.0130 0.0660 4.0430 0.6910 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 1.2770 0.8400 1.3070 1.6060 ;
      RECT 4.0130 0.9390 4.0430 1.6060 ;
      RECT 3.7090 0.0660 3.7390 0.6370 ;
      RECT 1.2770 0.0660 1.3070 0.6370 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 1.8850 0.0660 1.9150 0.6910 ;
      RECT 3.2530 0.0660 3.2830 0.6910 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 2.9490 0.8920 2.9790 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 3.7090 0.8390 3.7390 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
    LAYER NWELL ;
      RECT -0.1150 1.5430 8.6340 1.7730 ;
      RECT -0.1150 0.6980 5.4260 1.5430 ;
      RECT 8.3590 0.6790 8.6340 1.5430 ;
      RECT -0.1150 0.6790 4.4840 0.6980 ;
      RECT 4.9110 0.6790 5.4260 0.6980 ;
      RECT 5.8880 0.4910 7.8990 1.0830 ;
    LAYER M1 ;
      RECT 1.0230 0.5130 1.1650 0.5630 ;
      RECT 1.1150 0.5630 1.1650 0.7130 ;
      RECT 1.0390 0.7130 1.1650 0.7630 ;
      RECT 1.0390 0.7630 1.0890 1.0330 ;
      RECT 2.9990 0.3880 3.6730 0.4380 ;
      RECT 3.6230 0.4380 3.6730 0.5630 ;
      RECT 3.6230 0.2970 3.6730 0.3880 ;
      RECT 3.4710 0.9670 3.6890 1.0170 ;
      RECT 3.4710 0.4380 3.5210 0.9670 ;
      RECT 3.4710 1.0170 3.5210 1.1200 ;
      RECT 3.4710 1.1700 3.5210 1.2700 ;
      RECT 2.9990 1.1200 3.5210 1.1700 ;
      RECT 2.3890 0.8580 2.5490 0.9080 ;
      RECT 2.3890 0.9080 2.4390 0.9680 ;
      RECT 1.8590 0.9680 2.4390 1.0180 ;
      RECT 1.3430 0.8540 2.2450 0.9040 ;
      RECT 1.3430 0.9040 1.3930 1.0590 ;
      RECT 1.3430 0.6130 1.3930 0.8540 ;
      RECT 1.3430 1.0590 1.7130 1.1090 ;
      RECT 1.3430 0.5630 1.5450 0.6130 ;
      RECT 1.3430 1.1090 1.3930 1.3370 ;
      RECT 1.4950 0.4070 1.5450 0.5630 ;
      RECT 1.3430 0.4130 1.3930 0.5630 ;
      RECT 4.7630 0.6320 5.2850 0.6820 ;
      RECT 4.1190 0.4500 4.1690 0.7290 ;
      RECT 4.1190 0.7290 4.4850 0.7790 ;
      RECT 4.4350 0.7790 4.4850 1.1790 ;
      RECT 4.7630 0.6820 4.8130 0.6960 ;
      RECT 4.7630 0.4500 4.8130 0.6320 ;
      RECT 3.7750 0.4000 4.8130 0.4500 ;
      RECT 3.7760 1.1790 4.4850 1.2290 ;
      RECT 3.7750 0.4500 3.8250 0.5630 ;
      RECT 3.7750 0.2970 3.8250 0.4000 ;
      RECT 3.7760 1.2290 3.8260 1.3530 ;
      RECT 1.4030 1.3890 1.9410 1.4390 ;
      RECT 3.3230 0.1880 3.9170 0.2380 ;
      RECT 3.3230 0.2380 3.3730 0.2880 ;
      RECT 2.6820 0.2880 3.3730 0.3380 ;
      RECT 2.2950 0.4550 2.3450 0.6130 ;
      RECT 1.8590 0.6130 2.3450 0.6630 ;
      RECT 2.6820 0.3380 2.7320 0.4050 ;
      RECT 2.2950 0.4050 2.7320 0.4550 ;
      RECT 0.7950 1.5240 2.0930 1.5740 ;
      RECT 1.1910 0.8130 1.2810 0.8630 ;
      RECT 1.1910 0.8630 1.2410 1.0830 ;
      RECT 1.2310 0.4620 1.2810 0.8130 ;
      RECT 0.4310 1.0830 1.2410 1.1330 ;
      RECT 1.1750 0.4120 1.2810 0.4620 ;
      RECT 1.1910 1.1330 1.2410 1.3540 ;
      RECT 0.4310 0.7980 0.4810 1.0830 ;
      RECT 0.4310 0.7480 0.5210 0.7980 ;
      RECT 0.4310 0.4350 0.5210 0.4850 ;
      RECT 0.4310 0.3720 0.4810 0.4350 ;
      RECT 0.4710 0.4850 0.5210 0.7480 ;
      RECT 5.3370 0.6130 5.5890 0.6630 ;
      RECT 4.5350 0.8090 4.5850 1.3010 ;
      RECT 4.5350 0.5500 4.5850 0.7590 ;
      RECT 4.3070 0.5000 4.5850 0.5500 ;
      RECT 4.3070 0.5500 4.3570 0.6790 ;
      RECT 4.8390 0.8090 4.8890 1.3010 ;
      RECT 5.3370 0.6630 5.3870 0.7590 ;
      RECT 4.5350 0.7590 5.3870 0.8090 ;
      RECT 5.5070 1.1990 6.8050 1.2490 ;
      RECT 3.6230 0.8670 3.7650 0.9170 ;
      RECT 3.6230 0.6630 3.6730 0.8670 ;
      RECT 3.6230 0.6130 4.0690 0.6630 ;
      RECT 3.9340 0.9670 4.0690 1.0170 ;
      RECT 3.9340 0.9160 3.9840 0.9670 ;
      RECT 3.8350 0.8660 3.9840 0.9160 ;
      RECT 2.8470 0.4880 3.4080 0.5110 ;
      RECT 2.8470 0.5110 3.4090 0.5380 ;
      RECT 3.3590 0.5380 3.4090 1.0200 ;
      RECT 2.8630 1.0200 3.4090 1.0700 ;
      RECT 2.5990 0.7880 2.6490 1.1200 ;
      RECT 1.5500 0.7380 2.6510 0.7880 ;
      RECT 2.4070 0.5050 2.4570 0.7380 ;
      RECT 2.8630 1.0700 2.9130 1.1200 ;
      RECT 2.0870 1.1200 2.9130 1.1700 ;
      RECT 0.5830 0.6130 1.0290 0.6630 ;
      RECT 0.5830 0.6630 0.6330 1.0040 ;
      RECT 0.5830 0.4130 0.6330 0.6130 ;
      RECT 6.4950 0.8200 7.0430 0.8700 ;
      RECT 6.7990 0.7090 7.3370 0.7590 ;
      RECT 7.4230 0.6770 7.4730 0.7680 ;
      RECT 7.3830 0.4270 7.4730 0.4620 ;
      RECT 7.4230 0.1260 7.4730 0.4270 ;
      RECT 7.3830 0.6270 7.4730 0.6770 ;
      RECT 7.3830 0.5120 7.4330 0.6270 ;
      RECT 7.1790 0.4770 7.4330 0.5120 ;
      RECT 7.1790 0.4620 7.4730 0.4770 ;
      RECT 6.7990 0.1320 7.0330 0.1820 ;
      RECT 6.0550 1.0620 6.5040 1.1120 ;
      RECT 6.0550 0.6770 6.1050 1.0620 ;
      RECT 6.0150 0.6270 6.1050 0.6770 ;
      RECT 6.0150 0.4770 6.0650 0.6270 ;
      RECT 6.0150 0.4270 6.1050 0.4770 ;
      RECT 6.0550 0.1260 6.1050 0.4270 ;
      RECT 6.1150 0.5270 6.7130 0.5770 ;
      RECT 6.3590 0.5770 6.4090 0.8840 ;
      RECT 6.3590 0.1260 6.4090 0.5270 ;
      RECT 6.6630 0.5770 6.7130 0.7700 ;
      RECT 6.6630 0.3480 6.7130 0.5270 ;
      RECT 7.0270 1.0620 7.5650 1.1120 ;
      RECT 6.4950 0.2480 7.3370 0.2980 ;
      RECT 3.3770 1.5200 6.5010 1.5700 ;
      RECT 1.0980 0.0940 1.4910 0.1440 ;
      RECT 2.6190 1.5200 3.3090 1.5700 ;
      RECT 3.0740 0.6130 3.3090 0.6630 ;
      RECT 2.7110 0.9200 3.1410 0.9700 ;
      RECT 3.0910 0.8310 3.1410 0.9200 ;
      RECT 2.7110 0.9700 2.7610 1.0340 ;
      RECT 2.7110 0.5050 2.7610 0.9200 ;
      RECT 2.4670 1.4200 3.7730 1.4700 ;
      RECT 1.4790 1.1900 1.8650 1.2400 ;
      RECT 4.0560 1.2870 4.4490 1.3370 ;
  END
END RDFFNSRASRNX2_LVT

MACRO RDFFNSRASRQX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.36 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 8.3600 1.7020 ;
        RECT 0.2790 1.1310 0.3290 1.6420 ;
        RECT 2.1430 1.2700 2.1930 1.6420 ;
        RECT 0.4310 1.2940 0.4810 1.6420 ;
        RECT 6.3990 1.4540 6.4490 1.6420 ;
        RECT 1.9340 1.2200 3.2330 1.2700 ;
        RECT 0.4310 1.2440 0.9530 1.2940 ;
        RECT 3.9270 1.4040 6.4490 1.4540 ;
        RECT 3.9270 1.2790 3.9770 1.4040 ;
        RECT 4.9910 0.9590 5.0410 1.4040 ;
        RECT 4.6870 0.9530 4.7370 1.4040 ;
    END
  END VDD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.1430 0.9690 5.6770 1.0190 ;
        RECT 5.6270 0.3510 5.6770 0.9690 ;
        RECT 5.1430 1.0190 5.3750 1.1290 ;
        RECT 5.1270 0.3010 5.6770 0.3510 ;
        RECT 5.1430 1.1290 5.1930 1.3270 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 8.3600 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.2690 ;
        RECT 4.9910 0.0300 5.0410 0.2410 ;
        RECT 6.9670 0.0300 7.0170 0.1980 ;
        RECT 7.4230 0.0300 7.4730 0.4260 ;
        RECT 6.0550 0.0300 6.1050 0.4260 ;
        RECT 4.8630 0.0300 4.9130 0.2880 ;
        RECT 0.2790 0.2690 2.1530 0.3190 ;
        RECT 3.9110 0.2880 4.9130 0.3350 ;
        RECT 1.9510 0.3190 2.0010 0.5570 ;
        RECT 0.7350 0.3190 0.7850 0.5570 ;
        RECT 0.8870 0.3190 0.9370 0.5570 ;
        RECT 2.1030 0.3190 2.1530 0.5330 ;
        RECT 0.2790 0.3190 0.3290 0.4050 ;
        RECT 2.1030 0.2440 2.1530 0.2690 ;
        RECT 3.9110 0.3350 4.8880 0.3380 ;
        RECT 2.1030 0.1940 3.2330 0.2440 ;
        RECT 2.5590 0.2440 2.6090 0.3490 ;
    END
  END VSS

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.1550 0.8570 4.3110 0.9750 ;
        RECT 4.1550 0.9750 4.2050 1.0790 ;
        RECT 3.6230 1.0790 4.2050 1.1290 ;
        RECT 3.6230 1.1290 3.6730 1.3200 ;
        RECT 2.3310 1.3200 3.6730 1.3700 ;
        RECT 2.3310 1.3700 2.3810 1.4550 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6150 0.0880 4.6860 0.1380 ;
        RECT 1.6150 0.1380 1.7940 0.2100 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.4650 0.7250 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.4210 0.6630 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.5420 0.2490 7.6570 0.3590 ;
        RECT 7.5560 0.3590 7.6060 0.5270 ;
        RECT 7.3310 0.5270 7.6060 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8330 0.7030 2.9890 0.7310 ;
        RECT 2.8330 0.7310 3.2930 0.7810 ;
        RECT 2.9390 0.5970 2.9890 0.7030 ;
        RECT 2.8330 0.7810 2.9890 0.8150 ;
        RECT 3.2430 0.7810 3.2930 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 6.0390 0.9420 7.6570 1.0020 ;
        RECT 7.5470 0.6900 7.6570 0.9420 ;
        RECT 7.4230 0.6270 7.4730 0.9420 ;
    END
  END VDDG
  OBS
    LAYER PO ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 1.8850 0.9390 1.9150 1.6060 ;
      RECT 5.3810 0.0670 5.4110 1.6050 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 3.2530 0.8390 3.2830 1.6060 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 4.0130 0.0660 4.0430 0.6910 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 1.2770 0.8400 1.3070 1.6060 ;
      RECT 4.0130 0.9390 4.0430 1.6060 ;
      RECT 3.7090 0.0660 3.7390 0.6370 ;
      RECT 1.2770 0.0660 1.3070 0.6370 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 1.8850 0.0660 1.9150 0.6910 ;
      RECT 3.2530 0.0660 3.2830 0.6910 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 2.9490 0.8920 2.9790 1.6060 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 3.7090 0.8390 3.7390 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 2.9490 0.0660 2.9790 0.6910 ;
    LAYER NWELL ;
      RECT 5.7360 0.4910 7.7470 1.0830 ;
      RECT -0.1150 1.5430 8.4820 1.7730 ;
      RECT -0.1150 0.6790 5.2740 1.5430 ;
      RECT 8.2070 0.6790 8.4820 1.5430 ;
    LAYER M1 ;
      RECT 3.6230 0.2970 3.6730 0.3940 ;
      RECT 2.9990 0.3940 3.6730 0.4440 ;
      RECT 3.6230 0.4440 3.6730 0.5630 ;
      RECT 3.4710 0.9670 3.6890 1.0170 ;
      RECT 3.4710 0.4440 3.5210 0.9670 ;
      RECT 3.4710 1.0170 3.5210 1.1200 ;
      RECT 3.4710 1.1700 3.5210 1.2700 ;
      RECT 2.9990 1.1200 3.5210 1.1700 ;
      RECT 2.3890 0.8580 2.5490 0.9080 ;
      RECT 2.3890 0.9080 2.4390 0.9680 ;
      RECT 1.8590 0.9680 2.4390 1.0180 ;
      RECT 1.3430 0.8540 2.2450 0.9040 ;
      RECT 1.3430 0.9040 1.3930 1.0590 ;
      RECT 1.3430 0.6130 1.3930 0.8540 ;
      RECT 1.3430 1.0590 1.7130 1.1090 ;
      RECT 1.3430 0.5630 1.5450 0.6130 ;
      RECT 1.3430 1.1090 1.3930 1.3370 ;
      RECT 1.4950 0.4070 1.5450 0.5630 ;
      RECT 1.3430 0.4130 1.3930 0.5630 ;
      RECT 3.7750 0.4000 4.8130 0.4500 ;
      RECT 4.7630 0.4500 4.8130 0.6820 ;
      RECT 4.1190 0.4500 4.1690 0.7290 ;
      RECT 4.1190 0.7290 4.4850 0.7790 ;
      RECT 4.4350 0.7790 4.4850 1.1790 ;
      RECT 3.7760 1.1790 4.4850 1.2290 ;
      RECT 3.7750 0.4500 3.8250 0.5630 ;
      RECT 3.7750 0.2970 3.8250 0.4000 ;
      RECT 3.7760 1.2290 3.8260 1.3530 ;
      RECT 3.3230 0.1880 3.9170 0.2380 ;
      RECT 3.3230 0.2380 3.3730 0.2940 ;
      RECT 2.6820 0.2940 3.3730 0.3440 ;
      RECT 2.2950 0.4550 2.3450 0.6130 ;
      RECT 1.8590 0.6130 2.3450 0.6630 ;
      RECT 2.6820 0.3440 2.7320 0.4050 ;
      RECT 2.2950 0.4050 2.7320 0.4550 ;
      RECT 0.7950 1.5240 2.0930 1.5740 ;
      RECT 1.1910 0.8130 1.2810 0.8630 ;
      RECT 1.1910 0.8630 1.2410 1.0830 ;
      RECT 1.2310 0.4620 1.2810 0.8130 ;
      RECT 0.4310 1.0830 1.2410 1.1330 ;
      RECT 1.1750 0.4120 1.2810 0.4620 ;
      RECT 1.1910 1.1330 1.2410 1.3540 ;
      RECT 0.4310 0.7980 0.4810 1.0830 ;
      RECT 0.4310 0.7480 0.5210 0.7980 ;
      RECT 0.4310 0.4350 0.5210 0.4850 ;
      RECT 0.4310 0.3720 0.4810 0.4350 ;
      RECT 0.4710 0.4850 0.5210 0.7480 ;
      RECT 5.0150 0.6130 5.4370 0.6630 ;
      RECT 5.0150 0.6630 5.0650 0.7590 ;
      RECT 4.5350 0.7590 5.0650 0.8090 ;
      RECT 4.5350 0.8090 4.5850 1.3010 ;
      RECT 4.5350 0.5500 4.5850 0.7590 ;
      RECT 4.3070 0.5000 4.5850 0.5500 ;
      RECT 4.3070 0.5500 4.3570 0.6790 ;
      RECT 4.8390 0.8090 4.8890 1.3010 ;
      RECT 5.3550 1.1990 6.6530 1.2490 ;
      RECT 3.6230 0.8670 3.7650 0.9170 ;
      RECT 3.6230 0.6630 3.6730 0.8670 ;
      RECT 3.6230 0.6130 4.0690 0.6630 ;
      RECT 3.9340 0.9670 4.0690 1.0170 ;
      RECT 3.9340 0.9160 3.9840 0.9670 ;
      RECT 3.8350 0.8660 3.9840 0.9160 ;
      RECT 2.8470 0.4940 3.4080 0.5170 ;
      RECT 2.8470 0.5170 3.4090 0.5440 ;
      RECT 3.3590 0.5440 3.4090 1.0200 ;
      RECT 2.8630 1.0200 3.4090 1.0700 ;
      RECT 2.5990 0.7880 2.6490 1.1200 ;
      RECT 1.5500 0.7380 2.6510 0.7880 ;
      RECT 2.4070 0.5050 2.4570 0.7380 ;
      RECT 2.8630 1.0700 2.9130 1.1200 ;
      RECT 2.0870 1.1200 2.9130 1.1700 ;
      RECT 0.5830 0.6130 1.0290 0.6630 ;
      RECT 0.5830 0.6630 0.6330 1.0040 ;
      RECT 0.5830 0.4130 0.6330 0.6130 ;
      RECT 6.3430 0.8200 6.8910 0.8700 ;
      RECT 6.6470 0.7090 7.1850 0.7590 ;
      RECT 7.2710 0.6770 7.3210 0.7680 ;
      RECT 7.2310 0.4270 7.3210 0.4620 ;
      RECT 7.2710 0.1260 7.3210 0.4270 ;
      RECT 7.2310 0.6270 7.3210 0.6770 ;
      RECT 7.2310 0.5120 7.2810 0.6270 ;
      RECT 7.0270 0.4770 7.2810 0.5120 ;
      RECT 7.0270 0.4620 7.3210 0.4770 ;
      RECT 6.6470 0.1320 6.8810 0.1820 ;
      RECT 5.9030 1.0620 6.3520 1.1120 ;
      RECT 5.9030 0.6770 5.9530 1.0620 ;
      RECT 5.8630 0.6270 5.9530 0.6770 ;
      RECT 5.8630 0.4770 5.9130 0.6270 ;
      RECT 5.8630 0.4270 5.9530 0.4770 ;
      RECT 5.9030 0.1260 5.9530 0.4270 ;
      RECT 5.9630 0.5270 6.5610 0.5770 ;
      RECT 6.2070 0.5770 6.2570 0.8840 ;
      RECT 6.2070 0.1260 6.2570 0.5270 ;
      RECT 6.5110 0.5770 6.5610 0.7700 ;
      RECT 6.5110 0.3480 6.5610 0.5270 ;
      RECT 6.8750 1.0620 7.4130 1.1120 ;
      RECT 6.3430 0.2480 7.1850 0.2980 ;
      RECT 3.3770 1.5200 6.3490 1.5700 ;
      RECT 1.0980 0.0940 1.4910 0.1440 ;
      RECT 2.6190 1.5200 3.3090 1.5700 ;
      RECT 3.0740 0.6130 3.3090 0.6630 ;
      RECT 2.7110 0.9200 3.1410 0.9700 ;
      RECT 3.0910 0.8310 3.1410 0.9200 ;
      RECT 2.7110 0.9700 2.7610 1.0340 ;
      RECT 2.7110 0.5050 2.7610 0.9200 ;
      RECT 2.4670 1.4200 3.7730 1.4700 ;
      RECT 1.4790 1.1900 1.8650 1.2400 ;
      RECT 4.0560 1.2870 4.4490 1.3370 ;
      RECT 1.4030 1.3890 1.9410 1.4390 ;
      RECT 1.0390 0.7130 1.1650 0.7630 ;
      RECT 1.0390 0.7630 1.0890 1.0330 ;
      RECT 1.1150 0.5630 1.1650 0.7130 ;
      RECT 1.0230 0.5130 1.1650 0.5630 ;
  END
END RDFFNSRASRQX1_LVT

MACRO RDFFNSRASRQX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.512 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 8.5120 1.7020 ;
        RECT 0.2790 1.1310 0.3290 1.6420 ;
        RECT 2.1430 1.2700 2.1930 1.6420 ;
        RECT 0.4310 1.2940 0.4810 1.6420 ;
        RECT 6.5510 1.4540 6.6010 1.6420 ;
        RECT 1.9340 1.2200 3.2330 1.2700 ;
        RECT 0.4310 1.2440 0.9530 1.2940 ;
        RECT 3.9270 1.4040 6.6010 1.4540 ;
        RECT 3.9270 1.2790 3.9770 1.4040 ;
        RECT 4.9910 0.9590 5.0410 1.4040 ;
        RECT 4.6870 0.9530 4.7370 1.4040 ;
        RECT 5.2950 1.0690 5.3450 1.4040 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 8.5120 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.2690 ;
        RECT 4.9910 0.0300 5.0410 0.2410 ;
        RECT 5.2950 0.0300 5.3450 0.2410 ;
        RECT 7.1190 0.0300 7.1690 0.1980 ;
        RECT 7.5750 0.0300 7.6250 0.4260 ;
        RECT 6.2070 0.0300 6.2570 0.4260 ;
        RECT 4.8630 0.0300 4.9130 0.2880 ;
        RECT 0.2790 0.2690 2.1530 0.3190 ;
        RECT 3.9110 0.2880 4.9130 0.3380 ;
        RECT 1.9510 0.3190 2.0010 0.5570 ;
        RECT 0.7350 0.3190 0.7850 0.5570 ;
        RECT 0.8870 0.3190 0.9370 0.5570 ;
        RECT 2.1030 0.3190 2.1530 0.5330 ;
        RECT 0.2790 0.3190 0.3290 0.4050 ;
        RECT 2.1030 0.2380 2.1530 0.2690 ;
        RECT 2.1030 0.1880 3.2330 0.2380 ;
        RECT 2.5590 0.2380 2.6090 0.3490 ;
    END
  END VSS

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.1550 0.8570 4.3110 0.9750 ;
        RECT 4.1550 0.9750 4.2050 1.0790 ;
        RECT 3.6230 1.0790 4.2050 1.1290 ;
        RECT 3.6230 1.1290 3.6730 1.3200 ;
        RECT 2.3310 1.3200 3.6730 1.3700 ;
        RECT 2.3310 1.3700 2.3810 1.4550 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7230 0.0880 4.6610 0.0970 ;
        RECT 1.6150 0.0970 4.6610 0.1380 ;
        RECT 1.6150 0.1380 1.7730 0.2100 ;
        RECT 4.6110 0.1380 4.6610 0.1700 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.4650 0.7250 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.4210 0.6630 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.6950 0.2490 7.8090 0.3590 ;
        RECT 7.7080 0.3590 7.7580 0.5270 ;
        RECT 7.4830 0.5270 7.7580 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8330 0.7050 2.9890 0.7310 ;
        RECT 2.8330 0.7310 3.2930 0.7810 ;
        RECT 2.9390 0.5970 2.9890 0.7050 ;
        RECT 2.8330 0.7810 2.9890 0.8150 ;
        RECT 3.2430 0.7810 3.2930 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 6.1910 0.9420 7.8090 1.0020 ;
        RECT 7.6990 0.6900 7.8090 0.9420 ;
        RECT 7.5750 0.6270 7.6250 0.9420 ;
    END
  END VDDG

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.1430 0.9690 5.8290 1.0190 ;
        RECT 5.1430 1.0190 5.1930 1.3270 ;
        RECT 5.7790 0.3600 5.8290 0.9690 ;
        RECT 5.7190 0.3510 5.8330 0.3600 ;
        RECT 5.1270 0.3010 5.8330 0.3510 ;
        RECT 5.7190 0.2500 5.8330 0.3010 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q
  OBS
    LAYER PO ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 1.8850 0.9390 1.9150 1.6060 ;
      RECT 5.5330 0.0670 5.5630 1.6050 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 3.2530 0.8390 3.2830 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 4.0130 0.0660 4.0430 0.6910 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 1.2770 0.8400 1.3070 1.6060 ;
      RECT 4.0130 0.9390 4.0430 1.6060 ;
      RECT 3.7090 0.0660 3.7390 0.6370 ;
      RECT 1.2770 0.0660 1.3070 0.6370 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 1.8850 0.0660 1.9150 0.6910 ;
      RECT 3.2530 0.0660 3.2830 0.6910 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 2.9490 0.8920 2.9790 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 3.7090 0.8390 3.7390 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 2.9490 0.0660 2.9790 0.6910 ;
    LAYER NWELL ;
      RECT 5.8880 0.4910 7.8990 1.0830 ;
      RECT -0.1150 1.5430 8.6340 1.7730 ;
      RECT -0.1150 0.6790 5.4260 1.5430 ;
      RECT 8.3590 0.6790 8.6340 1.5430 ;
    LAYER M1 ;
      RECT 1.0390 0.7630 1.0890 1.0330 ;
      RECT 1.0390 0.7130 1.1650 0.7630 ;
      RECT 1.1150 0.5630 1.1650 0.7130 ;
      RECT 1.0230 0.5130 1.1650 0.5630 ;
      RECT 2.9990 0.3880 3.6730 0.4380 ;
      RECT 3.6230 0.4380 3.6730 0.5630 ;
      RECT 3.6230 0.2970 3.6730 0.3880 ;
      RECT 3.4710 0.9670 3.6890 1.0170 ;
      RECT 3.4710 0.4380 3.5210 0.9670 ;
      RECT 3.4710 1.0170 3.5210 1.1200 ;
      RECT 3.4710 1.1700 3.5210 1.2700 ;
      RECT 2.9990 1.1200 3.5210 1.1700 ;
      RECT 2.3890 0.8580 2.5490 0.9080 ;
      RECT 2.3890 0.9080 2.4390 0.9680 ;
      RECT 1.8590 0.9680 2.4390 1.0180 ;
      RECT 1.3430 0.8540 2.2450 0.9040 ;
      RECT 1.3430 0.9040 1.3930 1.0590 ;
      RECT 1.3430 0.6130 1.3930 0.8540 ;
      RECT 1.3430 1.0590 1.7130 1.1090 ;
      RECT 1.3430 0.5630 1.5450 0.6130 ;
      RECT 1.3430 1.1090 1.3930 1.3370 ;
      RECT 1.4950 0.4070 1.5450 0.5630 ;
      RECT 1.3430 0.4130 1.3930 0.5630 ;
      RECT 3.7750 0.4000 4.8130 0.4500 ;
      RECT 4.7630 0.4500 4.8130 0.6920 ;
      RECT 4.1190 0.4500 4.1690 0.7290 ;
      RECT 4.1190 0.7290 4.4850 0.7790 ;
      RECT 4.4350 0.7790 4.4850 1.1790 ;
      RECT 3.7760 1.1790 4.4850 1.2290 ;
      RECT 3.7750 0.4500 3.8250 0.5630 ;
      RECT 3.7750 0.2970 3.8250 0.4000 ;
      RECT 3.7760 1.2290 3.8260 1.3530 ;
      RECT 2.7110 0.9200 3.1410 0.9700 ;
      RECT 3.0910 0.8310 3.1410 0.9200 ;
      RECT 2.7110 0.9700 2.7610 1.0340 ;
      RECT 2.7110 0.5050 2.7610 0.9200 ;
      RECT 1.4790 1.1900 1.8650 1.2400 ;
      RECT 4.0560 1.2870 4.4490 1.3370 ;
      RECT 1.4030 1.3890 1.9410 1.4390 ;
      RECT 3.3230 0.1880 3.9170 0.2380 ;
      RECT 3.3230 0.2380 3.3730 0.2880 ;
      RECT 2.6820 0.2880 3.3730 0.3380 ;
      RECT 2.2950 0.4550 2.3450 0.6130 ;
      RECT 1.8590 0.6130 2.3450 0.6630 ;
      RECT 2.6820 0.3380 2.7320 0.4050 ;
      RECT 2.2950 0.4050 2.7320 0.4550 ;
      RECT 0.7950 1.5240 2.0930 1.5740 ;
      RECT 1.1910 0.8130 1.2810 0.8630 ;
      RECT 1.1910 0.8630 1.2410 1.0830 ;
      RECT 1.2310 0.4620 1.2810 0.8130 ;
      RECT 0.4310 1.0830 1.2410 1.1330 ;
      RECT 1.1750 0.4120 1.2810 0.4620 ;
      RECT 1.1910 1.1330 1.2410 1.3540 ;
      RECT 0.4310 0.7980 0.4810 1.0830 ;
      RECT 0.4310 0.7480 0.5210 0.7980 ;
      RECT 0.4310 0.4350 0.5210 0.4850 ;
      RECT 0.4310 0.3720 0.4810 0.4350 ;
      RECT 0.4710 0.4850 0.5210 0.7480 ;
      RECT 5.0150 0.6130 5.5890 0.6630 ;
      RECT 4.5350 0.8090 4.5850 1.3010 ;
      RECT 4.5350 0.5500 4.5850 0.7590 ;
      RECT 4.3070 0.5000 4.5850 0.5500 ;
      RECT 4.3070 0.5500 4.3570 0.6790 ;
      RECT 4.8390 0.8090 4.8890 1.3010 ;
      RECT 5.0150 0.6630 5.0650 0.7590 ;
      RECT 4.5350 0.7590 5.0650 0.8090 ;
      RECT 5.5070 1.1990 6.8050 1.2490 ;
      RECT 3.6230 0.8670 3.7650 0.9170 ;
      RECT 3.6230 0.6630 3.6730 0.8670 ;
      RECT 3.6230 0.6130 4.0690 0.6630 ;
      RECT 3.9340 0.9670 4.0690 1.0170 ;
      RECT 3.9340 0.9160 3.9840 0.9670 ;
      RECT 3.8350 0.8660 3.9840 0.9160 ;
      RECT 2.8470 0.4880 3.4090 0.5380 ;
      RECT 3.3590 0.5380 3.4090 1.0200 ;
      RECT 2.8630 1.0200 3.4090 1.0700 ;
      RECT 2.5990 0.7880 2.6490 1.1200 ;
      RECT 1.5500 0.7380 2.6510 0.7880 ;
      RECT 2.4070 0.5050 2.4570 0.7380 ;
      RECT 2.8630 1.0700 2.9130 1.1200 ;
      RECT 2.0870 1.1200 2.9130 1.1700 ;
      RECT 0.5830 0.6130 1.0290 0.6630 ;
      RECT 0.5830 0.6630 0.6330 1.0040 ;
      RECT 0.5830 0.4130 0.6330 0.6130 ;
      RECT 6.4950 0.8200 7.0430 0.8700 ;
      RECT 6.7990 0.7090 7.3370 0.7590 ;
      RECT 7.4230 0.6770 7.4730 0.7680 ;
      RECT 7.3830 0.4270 7.4730 0.4620 ;
      RECT 7.4230 0.1260 7.4730 0.4270 ;
      RECT 7.3830 0.6270 7.4730 0.6770 ;
      RECT 7.3830 0.5120 7.4330 0.6270 ;
      RECT 7.1790 0.4770 7.4330 0.5120 ;
      RECT 7.1790 0.4620 7.4730 0.4770 ;
      RECT 6.7990 0.1320 7.0330 0.1820 ;
      RECT 6.0550 1.0630 6.5040 1.1130 ;
      RECT 6.0550 0.6770 6.1050 1.0630 ;
      RECT 6.0150 0.6270 6.1050 0.6770 ;
      RECT 6.0150 0.4770 6.0650 0.6270 ;
      RECT 6.0150 0.4270 6.1050 0.4770 ;
      RECT 6.0550 0.1260 6.1050 0.4270 ;
      RECT 6.1150 0.5270 6.7130 0.5770 ;
      RECT 6.3590 0.5770 6.4090 0.8850 ;
      RECT 6.3590 0.1260 6.4090 0.5270 ;
      RECT 6.6630 0.5770 6.7130 0.7700 ;
      RECT 6.6630 0.3480 6.7130 0.5270 ;
      RECT 7.0270 1.0610 7.5650 1.1110 ;
      RECT 6.4950 0.2480 7.3370 0.2980 ;
      RECT 3.3770 1.5200 6.5010 1.5700 ;
      RECT 1.0980 0.0940 1.4910 0.1440 ;
      RECT 2.6190 1.5200 3.3090 1.5700 ;
      RECT 3.0740 0.6130 3.3090 0.6630 ;
      RECT 2.4670 1.4200 3.7730 1.4700 ;
  END
END RDFFNSRASRQX2_LVT

MACRO RDFFNSRASRX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.512 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 8.5120 1.7020 ;
        RECT 0.2790 1.1310 0.3290 1.6420 ;
        RECT 0.4480 1.2940 0.4980 1.6420 ;
        RECT 2.1430 1.2700 2.1930 1.6420 ;
        RECT 6.5510 1.4540 6.6010 1.6420 ;
        RECT 0.4480 1.2440 0.9530 1.2940 ;
        RECT 1.9340 1.2200 3.2330 1.2700 ;
        RECT 3.9270 1.4040 6.6010 1.4540 ;
        RECT 3.9270 1.2790 3.9770 1.4040 ;
        RECT 5.1430 0.9590 5.1930 1.4040 ;
        RECT 4.6870 0.9530 4.7370 1.4040 ;
    END
  END VDD

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.9910 0.4010 5.6910 0.4510 ;
        RECT 4.9910 0.1570 5.0410 0.4010 ;
        RECT 5.5690 0.4510 5.6910 0.5380 ;
        RECT 5.6410 0.5380 5.6910 0.8590 ;
        RECT 4.9910 0.8590 5.6910 0.9090 ;
        RECT 4.9910 0.9090 5.0410 1.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.2950 0.9690 5.8290 1.0190 ;
        RECT 5.7790 0.3510 5.8290 0.9690 ;
        RECT 5.2950 1.0190 5.5270 1.1290 ;
        RECT 5.2790 0.3010 5.8290 0.3510 ;
        RECT 5.2950 1.1290 5.3450 1.3270 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 8.5120 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.2640 ;
        RECT 5.1430 0.0300 5.1930 0.2410 ;
        RECT 7.1190 0.0300 7.1690 0.1980 ;
        RECT 7.5750 0.0300 7.6250 0.4260 ;
        RECT 6.2070 0.0300 6.2570 0.4260 ;
        RECT 4.8630 0.0300 4.9130 0.2880 ;
        RECT 0.2790 0.2640 2.1530 0.3140 ;
        RECT 3.9110 0.2880 4.9130 0.3380 ;
        RECT 1.9510 0.3140 2.0010 0.5570 ;
        RECT 0.7350 0.3140 0.7850 0.5570 ;
        RECT 0.8870 0.3140 0.9370 0.5570 ;
        RECT 2.1030 0.3140 2.1530 0.5330 ;
        RECT 0.2790 0.3140 0.3290 0.4050 ;
        RECT 2.1030 0.2380 2.1530 0.2640 ;
        RECT 2.1030 0.1880 3.2330 0.2380 ;
        RECT 2.5590 0.2380 2.6090 0.3490 ;
    END
  END VSS

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.1550 0.8570 4.3110 0.9750 ;
        RECT 4.1550 0.9750 4.2050 1.0790 ;
        RECT 3.6230 1.0790 4.2050 1.1290 ;
        RECT 3.6230 1.1290 3.6730 1.3200 ;
        RECT 2.3310 1.3200 3.6730 1.3700 ;
        RECT 2.3310 1.3700 2.3810 1.4550 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6150 0.0880 4.6610 0.1380 ;
        RECT 1.6150 0.1380 1.7730 0.2100 ;
        RECT 4.6110 0.1380 4.6610 0.1700 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.4210 0.6630 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN SAVE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.6940 0.2490 7.8090 0.3590 ;
        RECT 7.7080 0.3590 7.7580 0.5270 ;
        RECT 7.4830 0.5270 7.7580 0.5770 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SAVE

  PIN NRESTORE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8330 0.7040 2.9890 0.7310 ;
        RECT 2.8330 0.7310 3.2930 0.7810 ;
        RECT 2.9390 0.5970 2.9890 0.7040 ;
        RECT 2.8330 0.7810 2.9890 0.8150 ;
        RECT 3.2430 0.7810 3.2930 0.9330 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END NRESTORE

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.4650 0.7250 1.5750 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 6.1910 0.9420 7.8090 1.0020 ;
        RECT 7.6990 0.6900 7.8090 0.9420 ;
        RECT 7.5750 0.6270 7.6250 0.9420 ;
    END
  END VDDG
  OBS
    LAYER PO ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 7.0530 0.0660 7.0830 1.6060 ;
      RECT 2.9490 0.0660 2.9790 0.6910 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 1.8850 0.9390 1.9150 1.6060 ;
      RECT 5.5330 0.0670 5.5630 1.6050 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 7.2050 0.0660 7.2350 1.6060 ;
      RECT 5.9890 0.0660 6.0190 1.6060 ;
      RECT 3.2530 0.8390 3.2830 1.6060 ;
      RECT 7.6610 0.0660 7.6910 1.6060 ;
      RECT 6.9010 0.0660 6.9310 1.6060 ;
      RECT 7.3570 0.0660 7.3870 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 6.5970 0.0660 6.6270 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 4.0130 0.0660 4.0430 0.6910 ;
      RECT 6.2930 0.0660 6.3230 1.6060 ;
      RECT 1.5810 0.0660 1.6110 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 4.3170 0.0660 4.3470 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 1.7330 0.0660 1.7630 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 4.4690 0.0660 4.4990 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 1.2770 0.8400 1.3070 1.6060 ;
      RECT 4.0130 0.9390 4.0430 1.6060 ;
      RECT 3.7090 0.0660 3.7390 0.6370 ;
      RECT 1.2770 0.0660 1.3070 0.6370 ;
      RECT 7.5090 0.0660 7.5390 1.6060 ;
      RECT 1.8850 0.0660 1.9150 0.6910 ;
      RECT 3.2530 0.0660 3.2830 0.6910 ;
      RECT 6.1410 0.0660 6.1710 1.6060 ;
      RECT 7.8130 0.0660 7.8430 1.6060 ;
      RECT 2.9490 0.8920 2.9790 1.6060 ;
      RECT 6.4450 0.0660 6.4750 1.6060 ;
      RECT 5.8370 0.0660 5.8670 1.6060 ;
      RECT 3.7090 0.8390 3.7390 1.6060 ;
      RECT 7.9650 0.0660 7.9950 1.6060 ;
      RECT 8.4210 0.0660 8.4510 1.6060 ;
      RECT 6.7490 0.0660 6.7790 1.6060 ;
      RECT 8.1170 0.0660 8.1470 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 8.2690 0.0660 8.2990 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
    LAYER NWELL ;
      RECT 5.8880 0.4910 7.8990 1.0830 ;
      RECT -0.1150 1.5430 8.6340 1.7730 ;
      RECT -0.1150 0.6790 5.4260 1.5430 ;
      RECT 8.3590 0.6790 8.6340 1.5430 ;
    LAYER M1 ;
      RECT 1.0390 0.7130 1.1650 0.7630 ;
      RECT 1.0390 0.7630 1.0890 1.0330 ;
      RECT 1.1150 0.5630 1.1650 0.7130 ;
      RECT 1.0230 0.5130 1.1650 0.5630 ;
      RECT 2.9990 0.3880 3.6730 0.4380 ;
      RECT 3.6230 0.4380 3.6730 0.5630 ;
      RECT 3.6230 0.2970 3.6730 0.3880 ;
      RECT 3.4710 0.9670 3.6890 1.0170 ;
      RECT 3.4710 0.4380 3.5210 0.9670 ;
      RECT 3.4710 1.0170 3.5210 1.1200 ;
      RECT 3.4710 1.1700 3.5210 1.2700 ;
      RECT 2.9990 1.1200 3.5210 1.1700 ;
      RECT 2.3890 0.8580 2.5490 0.9080 ;
      RECT 2.3890 0.9080 2.4390 0.9680 ;
      RECT 1.8590 0.9680 2.4390 1.0180 ;
      RECT 1.3430 0.8540 2.2450 0.9040 ;
      RECT 1.3430 0.9040 1.3930 1.0590 ;
      RECT 1.3430 0.6130 1.3930 0.8540 ;
      RECT 1.3430 1.0590 1.7130 1.1090 ;
      RECT 1.3430 0.5630 1.5450 0.6130 ;
      RECT 1.3430 1.1090 1.3930 1.3370 ;
      RECT 1.4950 0.4070 1.5450 0.5630 ;
      RECT 1.3430 0.4130 1.3930 0.5630 ;
      RECT 4.7470 0.6320 5.1170 0.6820 ;
      RECT 5.0670 0.5970 5.1170 0.6320 ;
      RECT 4.1190 0.4500 4.1690 0.7290 ;
      RECT 4.1190 0.7290 4.4850 0.7790 ;
      RECT 4.4350 0.7790 4.4850 1.1790 ;
      RECT 4.7630 0.4500 4.8130 0.6320 ;
      RECT 3.7750 0.4000 4.8130 0.4500 ;
      RECT 3.7760 1.1790 4.4850 1.2290 ;
      RECT 3.7750 0.4500 3.8250 0.5630 ;
      RECT 3.7750 0.2970 3.8250 0.4000 ;
      RECT 3.7760 1.2290 3.8260 1.3530 ;
      RECT 0.7950 1.5240 2.0930 1.5740 ;
      RECT 1.1910 0.8130 1.2810 0.8630 ;
      RECT 1.1910 0.8630 1.2410 1.0830 ;
      RECT 1.2310 0.4620 1.2810 0.8130 ;
      RECT 0.4310 1.0830 1.2410 1.1330 ;
      RECT 1.1750 0.4120 1.2810 0.4620 ;
      RECT 1.1910 1.1330 1.2410 1.3540 ;
      RECT 0.4310 0.7980 0.4810 1.0830 ;
      RECT 0.4310 0.7480 0.5210 0.7980 ;
      RECT 0.4310 0.4350 0.5210 0.4850 ;
      RECT 0.4310 0.3720 0.4810 0.4350 ;
      RECT 0.4710 0.4850 0.5210 0.7480 ;
      RECT 3.3230 0.1880 3.9170 0.2380 ;
      RECT 3.3230 0.2380 3.3730 0.2880 ;
      RECT 2.6820 0.2880 3.3730 0.3380 ;
      RECT 2.2950 0.4550 2.3450 0.6130 ;
      RECT 1.8590 0.6130 2.3450 0.6630 ;
      RECT 2.6820 0.3380 2.7320 0.4050 ;
      RECT 2.2950 0.4050 2.7320 0.4550 ;
      RECT 5.1670 0.6130 5.5890 0.6630 ;
      RECT 4.5350 0.8090 4.5850 1.3010 ;
      RECT 4.5350 0.5500 4.5850 0.7590 ;
      RECT 4.3070 0.5000 4.5850 0.5500 ;
      RECT 4.3070 0.5500 4.3570 0.6790 ;
      RECT 4.8390 0.8090 4.8890 1.3010 ;
      RECT 5.1670 0.6630 5.2170 0.7590 ;
      RECT 4.5350 0.7590 5.2170 0.8090 ;
      RECT 5.5070 1.1990 6.8050 1.2490 ;
      RECT 3.6230 0.8670 3.7650 0.9170 ;
      RECT 3.6230 0.6630 3.6730 0.8670 ;
      RECT 3.6230 0.6130 4.0690 0.6630 ;
      RECT 3.9340 0.9670 4.0690 1.0170 ;
      RECT 3.9340 0.9160 3.9840 0.9670 ;
      RECT 3.8350 0.8660 3.9840 0.9160 ;
      RECT 2.8470 0.4880 3.4080 0.5110 ;
      RECT 2.8470 0.5110 3.4090 0.5380 ;
      RECT 3.3590 0.5380 3.4090 1.0200 ;
      RECT 2.8630 1.0200 3.4090 1.0700 ;
      RECT 2.5990 0.7880 2.6490 1.1200 ;
      RECT 1.5500 0.7380 2.6510 0.7880 ;
      RECT 2.4070 0.5050 2.4570 0.7380 ;
      RECT 2.8630 1.0700 2.9130 1.1200 ;
      RECT 2.0870 1.1200 2.9130 1.1700 ;
      RECT 0.5830 0.6130 1.0290 0.6630 ;
      RECT 0.5830 0.6630 0.6330 1.0040 ;
      RECT 0.5830 0.4130 0.6330 0.6130 ;
      RECT 6.4950 0.8200 7.0430 0.8700 ;
      RECT 6.7990 0.7090 7.3370 0.7590 ;
      RECT 7.4230 0.6770 7.4730 0.7680 ;
      RECT 7.3830 0.4270 7.4730 0.4620 ;
      RECT 7.4230 0.1260 7.4730 0.4270 ;
      RECT 7.3830 0.6270 7.4730 0.6770 ;
      RECT 7.3830 0.5120 7.4330 0.6270 ;
      RECT 7.1790 0.4770 7.4330 0.5120 ;
      RECT 7.1790 0.4620 7.4730 0.4770 ;
      RECT 6.7990 0.1320 7.0330 0.1820 ;
      RECT 6.0550 1.0620 6.5040 1.1120 ;
      RECT 6.0550 0.6770 6.1050 1.0620 ;
      RECT 6.0150 0.6270 6.1050 0.6770 ;
      RECT 6.0150 0.4770 6.0650 0.6270 ;
      RECT 6.0150 0.4270 6.1050 0.4770 ;
      RECT 6.0550 0.1260 6.1050 0.4270 ;
      RECT 6.1150 0.5270 6.7130 0.5770 ;
      RECT 6.3590 0.5770 6.4090 0.8840 ;
      RECT 6.3590 0.1260 6.4090 0.5270 ;
      RECT 6.6630 0.5770 6.7130 0.7700 ;
      RECT 6.6630 0.3480 6.7130 0.5270 ;
      RECT 7.0270 1.0620 7.5660 1.1120 ;
      RECT 6.4950 0.2480 7.3370 0.2980 ;
      RECT 3.3770 1.5200 6.5010 1.5700 ;
      RECT 1.0980 0.0940 1.4910 0.1440 ;
      RECT 2.6190 1.5200 3.3090 1.5700 ;
      RECT 3.0740 0.6130 3.3090 0.6630 ;
      RECT 2.7110 0.9200 3.1410 0.9700 ;
      RECT 3.0910 0.8310 3.1410 0.9200 ;
      RECT 2.7110 0.9700 2.7610 1.0340 ;
      RECT 2.7110 0.5050 2.7610 0.9200 ;
      RECT 2.4670 1.4200 3.7730 1.4700 ;
      RECT 1.4790 1.1900 1.8650 1.2400 ;
      RECT 4.0560 1.2870 4.4490 1.3370 ;
      RECT 1.4030 1.3890 1.9410 1.4390 ;
  END
END RDFFNSRASRX1_LVT

MACRO OR2X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.216 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8870 0.5110 1.0430 0.5580 ;
        RECT 0.8870 0.5080 1.1190 0.5110 ;
        RECT 0.9930 0.5580 1.0430 0.8160 ;
        RECT 0.9930 0.4010 1.1190 0.5080 ;
        RECT 0.8870 0.1990 0.9370 0.5080 ;
        RECT 0.8870 0.8160 1.0430 0.8660 ;
        RECT 0.8870 0.8660 0.9370 1.5440 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.2160 1.7020 ;
        RECT 0.7350 1.0860 0.7850 1.6420 ;
        RECT 0.2790 1.0870 0.3290 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.2160 0.0300 ;
        RECT 0.7350 0.0300 0.7850 0.3930 ;
        RECT 0.4310 0.0300 0.4810 0.3990 ;
    END
  END VSS

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5020 0.6420 0.6630 0.8150 ;
    END
    ANTENNAGATEAREA 0.0303 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.8570 0.4050 0.9670 ;
        RECT 0.3550 0.6420 0.4050 0.8570 ;
    END
    ANTENNAGATEAREA 0.0303 ;
  END A1
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.3310 1.7730 ;
    LAYER M1 ;
      RECT 0.7420 0.6580 0.8890 0.7080 ;
      RECT 0.7260 0.4860 0.7760 0.9560 ;
      RECT 0.5820 0.9050 0.7320 0.9550 ;
      RECT 0.2780 0.4860 0.7330 0.5360 ;
      RECT 0.5830 0.8890 0.6330 1.5250 ;
      RECT 0.5830 0.2990 0.6330 0.5120 ;
      RECT 0.2790 0.2970 0.3290 0.5120 ;
    LAYER PO ;
      RECT 1.1250 0.0730 1.1550 1.6000 ;
      RECT 0.9730 0.0730 1.0030 1.6000 ;
      RECT 0.0610 0.0730 0.0910 1.6040 ;
      RECT 0.8210 0.0730 0.8510 1.6040 ;
      RECT 0.2130 0.0730 0.2430 1.6040 ;
      RECT 0.6690 0.0730 0.6990 1.6040 ;
      RECT 0.3650 0.0730 0.3950 1.6040 ;
      RECT 0.5170 0.0730 0.5470 1.6040 ;
  END
END OR2X1_LVT

MACRO OR2X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.368 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8870 0.5450 1.2710 0.5950 ;
        RECT 0.8870 0.2080 0.9370 0.5450 ;
        RECT 1.1070 0.5950 1.2710 0.6630 ;
        RECT 1.1070 0.6630 1.1570 0.8400 ;
        RECT 0.8870 0.8400 1.1570 0.8900 ;
        RECT 0.8870 0.7970 0.9370 0.8400 ;
        RECT 0.8870 0.8900 0.9370 1.5250 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Y

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5050 0.6420 0.6630 0.8150 ;
    END
    ANTENNAGATEAREA 0.0306 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.8570 0.4050 0.9670 ;
        RECT 0.3550 0.6440 0.4050 0.8570 ;
    END
    ANTENNAGATEAREA 0.0306 ;
  END A1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.3680 1.7020 ;
        RECT 1.0390 0.9960 1.0890 1.6420 ;
        RECT 0.7350 1.0870 0.7850 1.6420 ;
        RECT 0.2790 1.0870 0.3290 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.3680 0.0300 ;
        RECT 0.7350 0.0300 0.7850 0.3820 ;
        RECT 1.0390 0.0300 1.0890 0.4740 ;
        RECT 0.4310 0.0300 0.4810 0.3990 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.4830 1.7730 ;
    LAYER M1 ;
      RECT 0.7810 0.6600 1.0290 0.7100 ;
      RECT 0.2790 0.3190 0.3290 0.5340 ;
      RECT 0.5830 0.9330 0.6330 1.5250 ;
      RECT 0.5830 0.3210 0.6330 0.5340 ;
      RECT 0.7560 0.5110 0.8060 0.9610 ;
      RECT 0.5830 0.9330 0.8060 0.9830 ;
      RECT 0.2780 0.4860 0.8060 0.5360 ;
    LAYER PO ;
      RECT 1.1250 0.0930 1.1550 1.6060 ;
      RECT 0.9730 0.0930 1.0030 1.6060 ;
      RECT 0.8210 0.0930 0.8510 1.6060 ;
      RECT 1.2770 0.0930 1.3070 1.6060 ;
      RECT 0.0610 0.0930 0.0910 1.6060 ;
      RECT 0.2130 0.0930 0.2430 1.6060 ;
      RECT 0.6690 0.0930 0.6990 1.6060 ;
      RECT 0.3650 0.0930 0.3950 1.6060 ;
      RECT 0.5170 0.0930 0.5470 1.6060 ;
  END
END OR2X2_LVT

MACRO OR2X4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.672 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8870 0.7970 0.9370 0.8210 ;
        RECT 0.8870 0.8210 1.4530 0.8710 ;
        RECT 0.8870 0.8710 0.9370 1.5400 ;
        RECT 1.1910 0.8710 1.2410 1.5400 ;
        RECT 1.1910 0.7970 1.2410 0.8210 ;
        RECT 1.4030 0.6630 1.4530 0.8210 ;
        RECT 1.4030 0.5950 1.5750 0.6630 ;
        RECT 0.8870 0.5530 1.5750 0.5950 ;
        RECT 0.8870 0.5450 1.4610 0.5530 ;
        RECT 0.8870 0.2080 0.9370 0.5450 ;
        RECT 1.1910 0.2080 1.2410 0.5450 ;
    END
    ANTENNADIFFAREA 0.2976 ;
  END Y

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5030 0.6310 0.6640 0.8150 ;
    END
    ANTENNAGATEAREA 0.0306 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2340 0.8570 0.4060 0.9670 ;
        RECT 0.3550 0.6220 0.4050 0.8570 ;
    END
    ANTENNAGATEAREA 0.0306 ;
  END A1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.6720 1.7020 ;
        RECT 1.3430 0.9680 1.3930 1.6420 ;
        RECT 1.0390 0.9680 1.0890 1.6420 ;
        RECT 0.7350 1.0490 0.7850 1.6420 ;
        RECT 0.2790 1.0700 0.3290 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.6720 0.0300 ;
        RECT 0.7350 0.0300 0.7850 0.3820 ;
        RECT 1.3430 0.0300 1.3930 0.4740 ;
        RECT 1.0390 0.0300 1.0890 0.4740 ;
        RECT 0.4310 0.0300 0.4810 0.3990 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.7870 1.7730 ;
    LAYER M1 ;
      RECT 0.7500 0.6580 1.3330 0.7080 ;
      RECT 0.2790 0.3190 0.3290 0.5340 ;
      RECT 0.5830 0.9330 0.6330 1.5250 ;
      RECT 0.5830 0.3210 0.6330 0.5340 ;
      RECT 0.7250 0.5110 0.7750 0.9610 ;
      RECT 0.5830 0.9330 0.7750 0.9830 ;
      RECT 0.2780 0.4860 0.7750 0.5360 ;
    LAYER PO ;
      RECT 1.2770 0.0930 1.3070 1.6040 ;
      RECT 1.4290 0.0930 1.4590 1.6040 ;
      RECT 1.1250 0.0930 1.1550 1.6040 ;
      RECT 0.9730 0.0930 1.0030 1.6040 ;
      RECT 0.8210 0.0930 0.8510 1.6040 ;
      RECT 0.0610 0.0930 0.0910 1.6040 ;
      RECT 1.5810 0.0930 1.6110 1.6040 ;
      RECT 0.2130 0.0930 0.2430 1.6040 ;
      RECT 0.6690 0.0930 0.6990 1.6040 ;
      RECT 0.3650 0.0930 0.3950 1.6040 ;
      RECT 0.5170 0.0930 0.5470 1.6040 ;
  END
END OR2X4_LVT

MACRO OR3X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.368 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 0.2490 1.2710 0.3590 ;
        RECT 1.1940 0.3590 1.2440 0.4260 ;
        RECT 1.0390 0.4260 1.2440 0.4760 ;
        RECT 1.0390 0.1310 1.0890 0.4260 ;
        RECT 1.0390 0.4760 1.0890 0.4920 ;
        RECT 1.1940 0.4760 1.2440 0.8030 ;
        RECT 1.0390 0.8030 1.2440 0.8530 ;
        RECT 1.0390 0.8530 1.0890 1.5340 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6600 0.5480 0.8150 0.7240 ;
    END
    ANTENNAGATEAREA 0.0285 ;
  END A3

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7050 0.4050 0.8150 ;
        RECT 0.3550 0.6420 0.4050 0.7050 ;
    END
    ANTENNAGATEAREA 0.0285 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5070 0.8570 0.6630 0.9670 ;
        RECT 0.5070 0.6420 0.5570 0.8570 ;
    END
    ANTENNAGATEAREA 0.0285 ;
  END A2

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.3680 1.7020 ;
        RECT 0.8870 0.9120 0.9370 1.6420 ;
        RECT 0.2790 0.9110 0.3290 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.3680 0.0300 ;
        RECT 0.8870 0.0300 0.9370 0.2950 ;
        RECT 0.7350 0.0300 0.7850 0.3240 ;
        RECT 0.4310 0.0300 0.4810 0.3240 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.4830 1.7730 ;
    LAYER M1 ;
      RECT 0.9010 0.6580 1.0290 0.7080 ;
      RECT 0.8810 0.3990 0.9310 0.8520 ;
      RECT 0.7350 0.8020 0.9060 0.8520 ;
      RECT 0.2790 0.3740 0.9310 0.4240 ;
      RECT 0.2790 0.3170 0.3290 0.3990 ;
      RECT 0.5830 0.3170 0.6330 0.3990 ;
      RECT 0.7350 0.8180 0.7850 1.5490 ;
    LAYER PO ;
      RECT 0.9730 0.0710 1.0030 1.6090 ;
      RECT 1.1250 0.0710 1.1550 1.6090 ;
      RECT 1.2770 0.0710 1.3070 1.6090 ;
      RECT 0.0610 0.0710 0.0910 1.6090 ;
      RECT 0.8210 0.0710 0.8510 1.6090 ;
      RECT 0.2130 0.0710 0.2430 1.6090 ;
      RECT 0.6690 0.0710 0.6990 1.6090 ;
      RECT 0.3650 0.0710 0.3950 1.6090 ;
      RECT 0.5170 0.0710 0.5470 1.6090 ;
  END
END OR3X1_LVT

MACRO OR3X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.52 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.5200 1.7020 ;
        RECT 1.1910 1.0040 1.2410 1.6420 ;
        RECT 0.8870 1.0040 0.9370 1.6420 ;
        RECT 0.2790 0.9110 0.3290 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.5200 0.0300 ;
        RECT 1.1910 0.0300 1.2410 0.3870 ;
        RECT 0.8870 0.0300 0.9370 0.2950 ;
        RECT 0.7350 0.0300 0.7850 0.3340 ;
        RECT 0.4310 0.0300 0.4810 0.3340 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6790 0.4050 0.8150 ;
        RECT 0.3550 0.6200 0.4050 0.6790 ;
    END
    ANTENNAGATEAREA 0.0285 ;
  END A1

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6600 0.5370 0.8150 0.7130 ;
    END
    ANTENNAGATEAREA 0.0285 ;
  END A3

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3130 0.4000 1.4230 0.4020 ;
        RECT 1.3030 0.4020 1.4230 0.5110 ;
        RECT 1.3030 0.5110 1.3530 0.5200 ;
        RECT 1.0390 0.5200 1.3530 0.5700 ;
        RECT 1.0390 0.1310 1.0890 0.5200 ;
        RECT 1.3030 0.5700 1.3530 0.8150 ;
        RECT 1.0390 0.8150 1.3530 0.8650 ;
        RECT 1.0390 0.8650 1.0890 1.5340 ;
        RECT 1.0390 0.8030 1.0890 0.8150 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Y

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5070 0.6300 0.5570 0.8570 ;
        RECT 0.5070 0.8570 0.6630 0.9670 ;
    END
    ANTENNAGATEAREA 0.0285 ;
  END A2
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.6350 1.7810 ;
    LAYER M1 ;
      RECT 0.8930 0.6560 1.1810 0.7060 ;
      RECT 0.5830 0.3290 0.6330 0.4110 ;
      RECT 0.7350 0.8170 0.7850 1.5480 ;
      RECT 0.8860 0.4110 0.9360 0.8800 ;
      RECT 0.2790 0.3860 0.9360 0.4360 ;
      RECT 0.7350 0.8300 0.9110 0.8800 ;
      RECT 0.2790 0.3290 0.3290 0.4110 ;
    LAYER PO ;
      RECT 1.4290 0.0920 1.4590 1.6210 ;
      RECT 0.9730 0.0710 1.0030 1.6210 ;
      RECT 1.1250 0.0710 1.1550 1.6210 ;
      RECT 1.2770 0.0920 1.3070 1.6210 ;
      RECT 0.0610 0.0920 0.0910 1.6210 ;
      RECT 0.8210 0.0920 0.8510 1.6210 ;
      RECT 0.2130 0.0920 0.2430 1.6210 ;
      RECT 0.6690 0.0920 0.6990 1.6210 ;
      RECT 0.3650 0.0920 0.3950 1.6210 ;
      RECT 0.5170 0.0920 0.5470 1.6210 ;
  END
END OR3X2_LVT

MACRO OR3X4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.432 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7050 0.4050 0.8150 ;
        RECT 0.3550 0.6450 0.4050 0.7050 ;
    END
    ANTENNAGATEAREA 0.0285 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5070 0.8570 0.6630 0.9670 ;
        RECT 0.5070 0.6450 0.5570 0.8570 ;
    END
    ANTENNAGATEAREA 0.0285 ;
  END A2

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.4320 1.7020 ;
        RECT 0.8870 0.9880 0.9370 1.6420 ;
        RECT 1.1910 0.9110 1.2410 1.6420 ;
        RECT 2.1030 1.0960 2.1530 1.6420 ;
        RECT 1.7990 1.0960 1.8490 1.6420 ;
        RECT 1.4950 1.0040 1.5450 1.6420 ;
        RECT 0.2790 0.9110 0.3290 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.4320 0.0300 ;
        RECT 2.1030 0.0300 2.1530 0.3870 ;
        RECT 1.4950 0.0300 1.5450 0.3870 ;
        RECT 0.8870 0.0300 0.9370 0.2030 ;
        RECT 1.1910 0.0300 1.2410 0.3870 ;
        RECT 1.7990 0.0300 1.8490 0.3870 ;
        RECT 0.7350 0.0300 0.7850 0.2440 ;
        RECT 0.4310 0.0300 0.4810 0.2440 ;
    END
  END VSS

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6600 0.5480 0.8150 0.7270 ;
    END
    ANTENNAGATEAREA 0.0285 ;
  END A3

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6310 0.9110 2.2850 0.9610 ;
        RECT 1.9510 0.9610 2.0010 1.5320 ;
        RECT 1.9510 0.8930 2.0010 0.9110 ;
        RECT 1.6470 0.9610 1.6970 1.5340 ;
        RECT 1.6470 0.8950 1.6970 0.9110 ;
        RECT 2.2340 0.5700 2.2840 0.9110 ;
        RECT 1.6470 0.5450 2.2840 0.5700 ;
        RECT 1.6470 0.5200 2.3350 0.5450 ;
        RECT 2.2250 0.4010 2.3350 0.5200 ;
        RECT 1.6470 0.1310 1.6970 0.5200 ;
        RECT 1.9510 0.1310 2.0010 0.5200 ;
    END
    ANTENNADIFFAREA 0.2976 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 2.5470 1.7730 ;
    LAYER M1 ;
      RECT 1.4970 0.6610 2.0930 0.7110 ;
      RECT 1.3430 0.1310 1.3930 0.5010 ;
      RECT 1.3430 0.8710 1.3930 1.5520 ;
      RECT 1.4970 0.5510 1.5470 0.6610 ;
      RECT 1.4970 0.7110 1.5470 0.8210 ;
      RECT 1.3430 0.5010 1.5470 0.5510 ;
      RECT 1.3430 0.8210 1.5470 0.8710 ;
      RECT 0.8770 0.6660 1.0290 0.7160 ;
      RECT 0.8770 0.3650 0.9270 0.6660 ;
      RECT 0.8770 0.7160 0.9270 0.8450 ;
      RECT 0.2790 0.3150 0.9270 0.3650 ;
      RECT 0.7350 0.8450 0.9270 0.8950 ;
      RECT 0.5830 0.2070 0.6330 0.3150 ;
      RECT 0.7350 0.8950 0.7850 1.5340 ;
      RECT 0.7350 0.8030 0.7850 0.8450 ;
      RECT 0.2790 0.2070 0.3290 0.3150 ;
      RECT 1.0390 0.5010 1.2120 0.5510 ;
      RECT 1.1620 0.5510 1.2120 0.6610 ;
      RECT 1.1620 0.6610 1.3330 0.7110 ;
      RECT 1.1620 0.7110 1.2120 0.7830 ;
      RECT 1.0390 0.7830 1.2120 0.8330 ;
      RECT 1.0390 0.1310 1.0890 0.5010 ;
      RECT 1.0390 0.8330 1.0890 1.1430 ;
    LAYER PO ;
      RECT 1.2770 0.0710 1.3070 1.6120 ;
      RECT 1.4290 0.0710 1.4590 1.6120 ;
      RECT 0.9730 0.0710 1.0030 1.6120 ;
      RECT 1.1250 0.0710 1.1550 1.6120 ;
      RECT 0.8210 0.0710 0.8510 1.6120 ;
      RECT 2.1890 0.0920 2.2190 1.6120 ;
      RECT 2.0370 0.0710 2.0670 1.6120 ;
      RECT 1.5810 0.0710 1.6110 1.6120 ;
      RECT 1.7330 0.0710 1.7630 1.6120 ;
      RECT 1.8850 0.0710 1.9150 1.6120 ;
      RECT 2.3410 0.0920 2.3710 1.6120 ;
      RECT 0.0610 0.0920 0.0910 1.6120 ;
      RECT 0.2130 0.0920 0.2430 1.6120 ;
      RECT 0.6690 0.0920 0.6990 1.6120 ;
      RECT 0.3650 0.0920 0.3950 1.6120 ;
      RECT 0.5170 0.0920 0.5470 1.6120 ;
  END
END OR3X4_LVT

MACRO OR4X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.128 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8110 0.6450 0.8610 0.7050 ;
        RECT 0.8110 0.7050 0.9670 0.8150 ;
    END
    ANTENNAGATEAREA 0.0279 ;
  END A4

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6590 0.4010 0.8150 0.5110 ;
        RECT 0.6590 0.5110 0.7090 0.7270 ;
    END
    ANTENNAGATEAREA 0.0279 ;
  END A3

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.1280 1.7020 ;
        RECT 1.0390 1.0650 1.0890 1.6420 ;
        RECT 1.3430 0.9110 1.3930 1.6420 ;
        RECT 1.6470 1.0960 1.6970 1.6420 ;
        RECT 0.2790 0.8130 0.3290 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.1280 0.0300 ;
        RECT 1.6470 0.0300 1.6970 0.3870 ;
        RECT 1.0390 0.0300 1.0890 0.2030 ;
        RECT 1.3430 0.0300 1.3930 0.3870 ;
        RECT 0.7350 0.0300 0.7850 0.2410 ;
        RECT 0.4310 0.0300 0.4810 0.2410 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6610 0.4210 0.7110 ;
        RECT 0.2490 0.5530 0.3590 0.6610 ;
    END
    ANTENNAGATEAREA 0.0279 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9190 0.2490 2.0310 0.3590 ;
        RECT 1.9190 0.3590 1.9690 0.4390 ;
        RECT 1.7990 0.4390 1.9690 0.4890 ;
        RECT 1.7990 0.1280 1.8490 0.4390 ;
        RECT 1.9190 0.4890 1.9690 0.7620 ;
        RECT 1.7990 0.7620 1.9690 0.8120 ;
        RECT 1.7990 0.8120 1.8490 1.5490 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5070 0.8570 0.6630 0.9670 ;
        RECT 0.5070 0.6450 0.5570 0.8570 ;
    END
    ANTENNAGATEAREA 0.0279 ;
  END A2
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 2.2430 1.8010 ;
    LAYER M1 ;
      RECT 1.0290 0.6660 1.1810 0.7160 ;
      RECT 1.0290 0.3410 1.0790 0.6660 ;
      RECT 1.0290 0.7160 1.0790 0.8980 ;
      RECT 0.8870 0.8980 1.0790 0.9480 ;
      RECT 0.2790 0.2910 1.0790 0.3410 ;
      RECT 0.5830 0.2100 0.6330 0.2910 ;
      RECT 0.8870 0.2090 0.9370 0.2910 ;
      RECT 0.8870 0.9480 0.9370 1.5500 ;
      RECT 0.2790 0.2100 0.3290 0.2910 ;
      RECT 1.3400 0.6610 1.4850 0.7110 ;
      RECT 1.3400 0.5520 1.3900 0.6610 ;
      RECT 1.3400 0.7110 1.3900 0.8030 ;
      RECT 1.1920 0.5270 1.3900 0.5520 ;
      RECT 1.1910 0.8030 1.3900 0.8530 ;
      RECT 1.1910 0.5020 1.3900 0.5270 ;
      RECT 1.1910 0.8530 1.2410 1.1520 ;
      RECT 1.1910 0.7920 1.2410 0.8030 ;
      RECT 1.1910 0.1310 1.2410 0.5020 ;
      RECT 1.6150 0.6610 1.7890 0.7110 ;
      RECT 1.4950 0.8970 1.6650 0.9470 ;
      RECT 1.6150 0.7110 1.6650 0.8970 ;
      RECT 1.6150 0.5520 1.6650 0.6610 ;
      RECT 1.4950 0.5020 1.6650 0.5520 ;
      RECT 1.4950 0.9470 1.5450 1.5350 ;
      RECT 1.4950 0.8810 1.5450 0.8970 ;
      RECT 1.4950 0.1280 1.5450 0.5020 ;
    LAYER PO ;
      RECT 1.1250 0.0710 1.1550 1.6120 ;
      RECT 1.2770 0.0710 1.3070 1.6120 ;
      RECT 1.4290 0.0710 1.4590 1.6100 ;
      RECT 1.5810 0.0720 1.6110 1.6100 ;
      RECT 0.9730 0.0720 1.0030 1.6100 ;
      RECT 0.0610 0.0720 0.0910 1.6100 ;
      RECT 2.0370 0.0720 2.0670 1.6100 ;
      RECT 0.8210 0.0720 0.8510 1.6100 ;
      RECT 1.8850 0.0720 1.9150 1.6100 ;
      RECT 1.7330 0.0710 1.7630 1.6100 ;
      RECT 0.2130 0.0720 0.2430 1.6100 ;
      RECT 0.6690 0.0720 0.6990 1.6100 ;
      RECT 0.3650 0.0720 0.3950 1.6100 ;
      RECT 0.5170 0.0720 0.5470 1.6100 ;
  END
END OR4X1_LVT

MACRO OR4X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.28 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0730 0.2490 2.1830 0.3590 ;
        RECT 2.1090 0.3590 2.1590 0.5030 ;
        RECT 1.7990 0.5030 2.1590 0.5530 ;
        RECT 1.7990 0.1310 1.8490 0.5030 ;
        RECT 2.1090 0.5530 2.1590 0.7880 ;
        RECT 1.7990 0.7880 2.1590 0.8380 ;
        RECT 1.7990 0.8380 1.8490 1.5520 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Y

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8090 0.7050 0.9670 0.8150 ;
        RECT 0.8110 0.6430 0.8610 0.7050 ;
    END
    ANTENNAGATEAREA 0.0279 ;
  END A4

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6590 0.4010 0.8150 0.5110 ;
        RECT 0.6590 0.5110 0.7090 0.7280 ;
    END
    ANTENNAGATEAREA 0.0279 ;
  END A3

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.2800 1.7020 ;
        RECT 1.9510 0.9110 2.0010 1.6420 ;
        RECT 1.6470 0.9120 1.6970 1.6420 ;
        RECT 1.0390 1.0650 1.0890 1.6420 ;
        RECT 1.3430 0.9120 1.3930 1.6420 ;
        RECT 0.2790 0.8180 0.3290 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.2800 0.0300 ;
        RECT 1.9510 0.0300 2.0010 0.3960 ;
        RECT 1.6470 0.0300 1.6970 0.3960 ;
        RECT 1.0390 0.0300 1.0890 0.2030 ;
        RECT 1.3430 0.0300 1.3930 0.3940 ;
        RECT 0.7350 0.0300 0.7850 0.2410 ;
        RECT 0.4310 0.0300 0.4810 0.2410 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6590 0.4210 0.7090 ;
        RECT 0.2490 0.5530 0.3590 0.6590 ;
    END
    ANTENNAGATEAREA 0.0279 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5070 0.8570 0.6630 0.9670 ;
        RECT 0.5070 0.6430 0.5570 0.8570 ;
    END
    ANTENNAGATEAREA 0.0279 ;
  END A2
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 2.3950 1.8010 ;
    LAYER M1 ;
      RECT 1.0290 0.6660 1.1810 0.7160 ;
      RECT 1.0290 0.3410 1.0790 0.6660 ;
      RECT 1.0290 0.7160 1.0790 0.9270 ;
      RECT 0.8870 0.9270 1.0790 0.9770 ;
      RECT 0.2790 0.2910 1.0790 0.3410 ;
      RECT 0.5830 0.2100 0.6330 0.2910 ;
      RECT 0.8870 0.2090 0.9370 0.2910 ;
      RECT 0.8870 0.9770 0.9370 1.5350 ;
      RECT 0.2790 0.2100 0.3290 0.2910 ;
      RECT 1.3400 0.6610 1.4850 0.7110 ;
      RECT 1.3400 0.5520 1.3900 0.6610 ;
      RECT 1.3400 0.7110 1.3900 0.8030 ;
      RECT 1.1910 0.5020 1.3900 0.5520 ;
      RECT 1.1910 0.8030 1.3900 0.8530 ;
      RECT 1.1910 0.1310 1.2410 0.5020 ;
      RECT 1.1910 0.8530 1.2410 1.0510 ;
      RECT 1.1910 0.7830 1.2410 0.8030 ;
      RECT 1.6180 0.6610 1.9410 0.7110 ;
      RECT 1.4950 0.1280 1.5450 0.5030 ;
      RECT 1.4950 0.8530 1.5450 1.5350 ;
      RECT 1.4950 0.7890 1.5450 0.8030 ;
      RECT 1.6180 0.5530 1.6680 0.6610 ;
      RECT 1.6180 0.7110 1.6680 0.8030 ;
      RECT 1.4950 0.5030 1.6680 0.5530 ;
      RECT 1.4950 0.8030 1.6680 0.8530 ;
    LAYER PO ;
      RECT 1.7330 0.0710 1.7630 1.6120 ;
      RECT 1.8850 0.0710 1.9150 1.6120 ;
      RECT 2.0370 0.0710 2.0670 1.6120 ;
      RECT 1.5810 0.0710 1.6110 1.6120 ;
      RECT 1.1250 0.0710 1.1550 1.6120 ;
      RECT 1.2770 0.0710 1.3070 1.6120 ;
      RECT 1.4290 0.0710 1.4590 1.6100 ;
      RECT 0.9730 0.0720 1.0030 1.6100 ;
      RECT 0.0610 0.0720 0.0910 1.6100 ;
      RECT 2.1890 0.0720 2.2190 1.6100 ;
      RECT 0.8210 0.0720 0.8510 1.6100 ;
      RECT 0.2130 0.0720 0.2430 1.6100 ;
      RECT 0.6690 0.0720 0.6990 1.6100 ;
      RECT 0.3650 0.0720 0.3950 1.6100 ;
      RECT 0.5170 0.0720 0.5470 1.6100 ;
  END
END OR4X2_LVT

MACRO OR4X4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.584 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3770 0.2490 2.4870 0.3590 ;
        RECT 2.3890 0.3590 2.4390 0.4400 ;
        RECT 1.7990 0.4400 2.4390 0.4900 ;
        RECT 2.1030 0.4900 2.1530 0.4920 ;
        RECT 2.1030 0.1310 2.1530 0.4400 ;
        RECT 1.7990 0.1310 1.8490 0.4400 ;
        RECT 1.7990 0.4900 1.8490 0.4920 ;
        RECT 2.3890 0.4900 2.4390 0.8950 ;
        RECT 1.7990 0.8950 2.4390 0.9450 ;
        RECT 2.1030 0.9450 2.1530 1.5340 ;
        RECT 1.7990 0.9450 1.8490 1.5340 ;
    END
    ANTENNADIFFAREA 0.2976 ;
  END Y

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8070 0.4000 0.9670 0.5110 ;
        RECT 0.8110 0.5110 0.8610 0.6070 ;
    END
    ANTENNAGATEAREA 0.0315 ;
  END A4

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6570 0.7050 0.8150 0.8150 ;
        RECT 0.6590 0.5250 0.7090 0.7050 ;
    END
    ANTENNAGATEAREA 0.0315 ;
  END A3

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.5840 1.7020 ;
        RECT 2.2550 1.0950 2.3050 1.6420 ;
        RECT 1.9510 1.0960 2.0010 1.6420 ;
        RECT 1.6470 1.0960 1.6970 1.6420 ;
        RECT 1.0390 0.8810 1.0890 1.6420 ;
        RECT 1.3430 1.0050 1.3930 1.6420 ;
        RECT 0.2790 0.7240 0.3290 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.5840 0.0300 ;
        RECT 1.3430 0.0300 1.3930 0.3190 ;
        RECT 2.2550 0.0300 2.3050 0.3180 ;
        RECT 1.6470 0.0300 1.6970 0.3190 ;
        RECT 1.9510 0.0300 2.0010 0.3190 ;
        RECT 1.0390 0.0300 1.0890 0.2030 ;
        RECT 0.7350 0.0300 0.7850 0.2000 ;
        RECT 0.4310 0.0300 0.4810 0.2000 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5250 0.4200 0.6630 ;
    END
    ANTENNAGATEAREA 0.0315 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 0.8570 0.5570 0.9670 ;
        RECT 0.5070 0.5250 0.5570 0.8570 ;
    END
    ANTENNAGATEAREA 0.0315 ;
  END A2
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 2.6990 1.8010 ;
      RECT 0.1980 0.5620 1.0180 0.6790 ;
    LAYER M1 ;
      RECT 1.6180 0.6610 2.2450 0.7110 ;
      RECT 1.4950 0.9470 1.5450 1.5350 ;
      RECT 1.4950 0.8810 1.5450 0.8970 ;
      RECT 1.4950 0.5560 1.5450 0.5570 ;
      RECT 1.4950 0.1280 1.5450 0.5060 ;
      RECT 1.6180 0.7110 1.6680 0.8970 ;
      RECT 1.6180 0.5560 1.6680 0.6610 ;
      RECT 1.4950 0.8970 1.6680 0.9470 ;
      RECT 1.4950 0.5060 1.6680 0.5560 ;
      RECT 1.0290 0.6660 1.1810 0.7160 ;
      RECT 1.0290 0.3030 1.0790 0.6660 ;
      RECT 1.0290 0.7160 1.0790 0.7310 ;
      RECT 0.8870 0.7310 1.0790 0.7810 ;
      RECT 0.2790 0.2530 1.0790 0.3030 ;
      RECT 0.5830 0.1690 0.6330 0.2530 ;
      RECT 0.8870 0.1680 0.9370 0.2530 ;
      RECT 0.8870 0.7810 0.9370 1.5350 ;
      RECT 0.2790 0.1690 0.3290 0.2530 ;
      RECT 1.3400 0.6610 1.4850 0.7110 ;
      RECT 1.3400 0.4770 1.3900 0.6610 ;
      RECT 1.3400 0.7110 1.3900 0.8030 ;
      RECT 1.1920 0.4520 1.3900 0.4770 ;
      RECT 1.1910 0.8030 1.3900 0.8530 ;
      RECT 1.1910 0.4270 1.3900 0.4520 ;
      RECT 1.1910 0.8530 1.2410 1.0510 ;
      RECT 1.1910 0.7830 1.2410 0.8030 ;
      RECT 1.1910 0.1310 1.2410 0.4270 ;
    LAYER PO ;
      RECT 2.0370 0.0710 2.0670 1.6120 ;
      RECT 1.8850 0.0710 1.9150 1.6120 ;
      RECT 1.7330 0.0710 1.7630 1.6120 ;
      RECT 2.1890 0.0710 2.2190 1.6120 ;
      RECT 2.3410 0.0710 2.3710 1.6120 ;
      RECT 1.5810 0.0710 1.6110 1.6120 ;
      RECT 1.1250 0.0710 1.1550 1.6120 ;
      RECT 1.2770 0.0710 1.3070 1.6120 ;
      RECT 1.4290 0.0710 1.4590 1.6100 ;
      RECT 0.9730 0.0610 1.0030 1.6100 ;
      RECT 0.0610 0.0610 0.0910 1.6100 ;
      RECT 2.4930 0.0720 2.5230 1.6100 ;
      RECT 0.8210 0.0610 0.8510 1.6100 ;
      RECT 0.2130 0.0610 0.2430 1.6100 ;
      RECT 0.6690 0.0610 0.6990 1.6100 ;
      RECT 0.3650 0.0610 0.3950 1.6100 ;
      RECT 0.5170 0.0610 0.5470 1.6100 ;
  END
END OR4X4_LVT

MACRO PGX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.76 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 0.7600 1.7020 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 0.7600 0.0300 ;
    END
  END VSS

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0970 0.0920 0.4360 0.1420 ;
        RECT 0.0970 0.1420 0.2070 0.2050 ;
    END
    ANTENNAGATEAREA 0.01125 ;
  END AN

  PIN INOUT1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0970 0.5530 0.3290 0.6630 ;
        RECT 0.2790 0.6630 0.3290 1.4720 ;
        RECT 0.2790 0.1920 0.3290 0.5530 ;
    END
    ANTENNADIFFAREA 0.1111 ;
    ANTENNAGATEAREA 0.1111 ;
  END INOUT1

  PIN INOUT2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4310 0.1920 0.4810 0.7050 ;
        RECT 0.4310 0.7050 0.6630 0.8150 ;
        RECT 0.4310 0.8150 0.4810 1.4720 ;
    END
    ANTENNADIFFAREA 0.1111 ;
    ANTENNAGATEAREA 0.1111 ;
  END INOUT2

  PIN AP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3240 1.5280 0.6630 1.5780 ;
        RECT 0.5530 1.4650 0.6630 1.5280 ;
    END
    ANTENNAGATEAREA 0.02145 ;
  END AP
  OBS
    LAYER NWELL ;
      RECT -0.1120 0.6790 0.8720 1.7730 ;
    LAYER PO ;
      RECT 0.3650 0.7170 0.3950 1.6060 ;
      RECT 0.3650 0.0640 0.3950 0.6150 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
  END
END PGX1_LVT

MACRO PGX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.912 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 0.9120 1.7020 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 0.9120 0.0300 ;
    END
  END VSS

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0970 0.0920 0.5880 0.1420 ;
        RECT 0.0970 0.1420 0.2070 0.2070 ;
    END
    ANTENNAGATEAREA 0.0225 ;
  END AN

  PIN INOUT1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0970 0.5530 0.3290 0.6630 ;
        RECT 0.2790 0.6630 0.3290 1.4280 ;
        RECT 0.2790 0.1920 0.3290 0.5530 ;
        RECT 0.2790 1.4280 0.6330 1.4780 ;
        RECT 0.5830 0.3080 0.6330 1.4280 ;
    END
    ANTENNADIFFAREA 0.2222 ;
    ANTENNAGATEAREA 0.2222 ;
  END INOUT1

  PIN INOUT2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4310 0.1920 0.7330 0.2420 ;
        RECT 0.6830 0.2420 0.7330 0.2490 ;
        RECT 0.4310 0.2420 0.4810 1.3780 ;
        RECT 0.6830 0.2490 0.8150 0.3590 ;
    END
    ANTENNADIFFAREA 0.133 ;
    ANTENNAGATEAREA 0.133 ;
  END INOUT2

  PIN AP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3240 1.5280 0.8150 1.5780 ;
        RECT 0.7050 1.4650 0.8150 1.5280 ;
    END
    ANTENNAGATEAREA 0.0429 ;
  END AP
  OBS
    LAYER NWELL ;
      RECT -0.1120 0.6790 1.0240 1.7730 ;
    LAYER PO ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
      RECT 0.5170 0.0660 0.5470 0.6150 ;
      RECT 0.5170 0.7170 0.5470 1.6060 ;
      RECT 0.3650 0.7170 0.3950 1.6060 ;
      RECT 0.3650 0.0640 0.3950 0.6150 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
  END
END PGX2_LVT

MACRO PGX4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.216 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.2160 1.7020 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.2160 0.0300 ;
    END
  END VSS

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0970 0.0920 0.8920 0.1420 ;
        RECT 0.0970 0.1420 0.2070 0.2070 ;
    END
    ANTENNAGATEAREA 0.045 ;
  END AN

  PIN INOUT1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0970 0.5530 0.3290 0.6630 ;
        RECT 0.2790 0.6630 0.3290 1.4280 ;
        RECT 0.2790 0.1920 0.3290 0.5530 ;
        RECT 0.2790 1.4280 0.9370 1.4780 ;
        RECT 0.8870 0.3080 0.9370 1.4280 ;
        RECT 0.5830 0.3080 0.6330 1.4280 ;
    END
    ANTENNADIFFAREA 0.3552 ;
    ANTENNAGATEAREA 0.3552 ;
  END INOUT1

  PIN INOUT2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4310 0.1920 1.0370 0.2420 ;
        RECT 0.9870 0.2420 1.0370 0.2490 ;
        RECT 0.7350 0.2420 0.7850 1.3780 ;
        RECT 0.4310 0.2420 0.4810 1.3780 ;
        RECT 0.9870 0.2490 1.1190 0.3590 ;
    END
    ANTENNADIFFAREA 0.266 ;
    ANTENNAGATEAREA 0.266 ;
  END INOUT2

  PIN AP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3240 1.5280 1.1190 1.5780 ;
        RECT 1.0090 1.4650 1.1190 1.5280 ;
    END
    ANTENNAGATEAREA 0.0858 ;
  END AP
  OBS
    LAYER NWELL ;
      RECT -0.1120 0.6790 1.3280 1.7730 ;
    LAYER PO ;
      RECT 0.6690 0.0660 0.6990 0.6150 ;
      RECT 0.6690 0.7170 0.6990 1.6060 ;
      RECT 0.8210 0.0660 0.8510 0.6150 ;
      RECT 0.8210 0.7170 0.8510 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 0.5170 0.0660 0.5470 0.6150 ;
      RECT 0.5170 0.7170 0.5470 1.6060 ;
      RECT 0.3650 0.7170 0.3950 1.6060 ;
      RECT 0.3650 0.0640 0.3950 0.6150 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
  END
END PGX4_LVT

MACRO PMT1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.76 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.8570 0.3590 0.9670 ;
        RECT 0.2790 0.9670 0.3290 1.5550 ;
        RECT 0.2790 0.8290 0.3290 0.8570 ;
    END
    ANTENNADIFFAREA 0.0816 ;
    ANTENNAGATEAREA 0.0816 ;
  END S

  PIN D
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 1.4590 0.5110 1.5750 ;
        RECT 0.4310 0.8290 0.4810 1.4590 ;
    END
    ANTENNADIFFAREA 0.0816 ;
  END D

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 0.7600 0.0300 ;
    END
  END VSS

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.6590 0.5110 0.7090 ;
        RECT 0.4010 0.5530 0.5110 0.6590 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END G

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 0.7600 1.7020 ;
    END
  END VDD
  OBS
    LAYER NWELL ;
      RECT -0.1250 0.6790 0.8650 1.7730 ;
    LAYER PO ;
      RECT 0.3650 0.6430 0.3950 1.6050 ;
      RECT 0.5170 0.6430 0.5470 1.6010 ;
      RECT 0.6690 0.6430 0.6990 1.6010 ;
      RECT 0.0610 0.6430 0.0910 1.6050 ;
      RECT 0.2130 0.6430 0.2430 1.6050 ;
  END
END PMT1_LVT

MACRO OA221X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.976 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.9760 0.0300 ;
        RECT 1.4950 0.0300 1.5450 0.3990 ;
        RECT 0.4310 0.0300 0.4810 0.5120 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7100 0.4210 0.8170 ;
        RECT 0.2490 0.7010 0.3590 0.7100 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END A1

  PIN A5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0230 0.5410 1.1230 0.5490 ;
        RECT 1.0090 0.5490 1.1230 0.6010 ;
        RECT 1.0090 0.6010 1.1650 0.6750 ;
        RECT 1.1150 0.6750 1.1650 0.8080 ;
    END
    ANTENNAGATEAREA 0.0177 ;
  END A5

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.9760 1.7020 ;
        RECT 0.8870 1.3350 0.9370 1.6420 ;
        RECT 1.0390 1.3330 1.0890 1.6420 ;
        RECT 1.4950 1.1330 1.5450 1.6420 ;
        RECT 0.2790 0.9580 0.3290 1.6420 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3430 0.5300 1.8360 0.5420 ;
        RECT 1.7860 0.5420 1.8360 0.9560 ;
        RECT 1.3430 0.4920 1.9110 0.5300 ;
        RECT 1.3430 0.9560 1.8360 1.0060 ;
        RECT 1.7510 0.3920 1.9110 0.4920 ;
        RECT 1.6470 0.1880 1.6970 0.4920 ;
        RECT 1.3430 0.1880 1.3930 0.4920 ;
        RECT 1.6470 1.0060 1.6970 1.4260 ;
        RECT 1.3430 1.0060 1.3930 1.4260 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END Y

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 1.4610 0.5730 1.5750 ;
        RECT 0.4260 1.4600 0.5730 1.4610 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8110 0.8420 0.8610 1.0020 ;
        RECT 0.8110 1.0020 0.9680 1.1390 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END A3

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6590 0.7130 0.7090 0.8540 ;
        RECT 0.5530 0.8540 0.7090 0.9860 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END A4
  OBS
    LAYER NWELL ;
      RECT -0.1350 0.6790 2.0920 1.7870 ;
    LAYER M1 ;
      RECT 1.5350 0.6810 1.6210 0.6990 ;
      RECT 1.2270 0.6310 1.6210 0.6810 ;
      RECT 1.5350 0.6130 1.6210 0.6310 ;
      RECT 1.2270 0.5330 1.2770 0.6310 ;
      RECT 1.2270 0.6810 1.2770 0.9030 ;
      RECT 1.1910 0.4830 1.2770 0.5330 ;
      RECT 1.0390 0.9030 1.2770 0.9530 ;
      RECT 1.1910 0.2110 1.2410 0.4830 ;
      RECT 1.1910 0.9530 1.2410 1.4270 ;
      RECT 1.0390 0.9530 1.0890 1.2130 ;
      RECT 0.5830 1.2130 1.0890 1.2630 ;
      RECT 1.3830 0.6810 1.4690 0.6990 ;
      RECT 1.3830 0.6130 1.4690 0.6310 ;
      RECT 0.5830 1.2630 0.6330 1.3930 ;
      RECT 0.5830 1.1060 0.6330 1.2130 ;
      RECT 0.7350 0.0980 1.0890 0.1480 ;
      RECT 1.0390 0.1480 1.0890 0.4310 ;
      RECT 0.7350 0.1480 0.7850 0.5010 ;
      RECT 0.2790 0.5980 0.9370 0.6480 ;
      RECT 0.5830 0.1810 0.6330 0.5980 ;
      RECT 0.8870 0.2080 0.9370 0.5980 ;
      RECT 0.2790 0.1780 0.3290 0.5980 ;
    LAYER PO ;
      RECT 1.1250 0.1010 1.1550 1.4690 ;
      RECT 1.8850 0.1010 1.9150 1.4690 ;
      RECT 0.5170 0.1010 0.5470 1.5670 ;
      RECT 1.5810 0.0690 1.6110 1.6080 ;
      RECT 0.8210 0.1010 0.8510 1.4690 ;
      RECT 0.6690 0.1010 0.6990 1.4690 ;
      RECT 0.2130 0.1010 0.2430 1.4690 ;
      RECT 0.3650 0.1010 0.3950 1.4690 ;
      RECT 1.2770 0.1010 1.3070 1.4690 ;
      RECT 1.7330 0.1010 1.7630 1.4690 ;
      RECT 1.4290 0.0690 1.4590 1.6080 ;
      RECT 0.9730 0.1010 1.0030 1.4690 ;
      RECT 0.0610 0.1010 0.0910 1.4690 ;
  END
END OA221X2_LVT

MACRO OA222X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.976 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6590 0.7130 0.7090 0.8540 ;
        RECT 0.5530 0.8540 0.7090 0.9860 ;
    END
    ANTENNAGATEAREA 0.0231 ;
  END A4

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8110 0.8420 0.8610 1.0020 ;
        RECT 0.8110 1.0020 0.9680 1.1390 ;
    END
    ANTENNAGATEAREA 0.0231 ;
  END A3

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 1.4610 0.5730 1.5750 ;
        RECT 0.4260 1.4600 0.5730 1.4610 ;
    END
    ANTENNAGATEAREA 0.0231 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7100 0.4210 0.8170 ;
        RECT 0.2490 0.7010 0.3590 0.7100 ;
    END
    ANTENNAGATEAREA 0.0231 ;
  END A1

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.9760 0.0300 ;
        RECT 0.4310 0.0300 0.4810 0.5120 ;
        RECT 1.4950 0.0300 1.5450 0.3990 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.9760 1.7020 ;
        RECT 1.4950 1.1330 1.5450 1.6420 ;
        RECT 1.0390 1.3330 1.0890 1.6420 ;
        RECT 0.2790 0.9580 0.3290 1.6420 ;
        RECT 0.8870 1.3350 0.9370 1.6420 ;
    END
  END VDD

  PIN A6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1600 1.1570 1.2800 1.2810 ;
        RECT 1.1710 1.1460 1.2800 1.1570 ;
        RECT 1.1710 1.2810 1.2210 1.4850 ;
        RECT 1.1710 1.4850 1.3390 1.5350 ;
    END
    ANTENNAGATEAREA 0.0231 ;
  END A6

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6470 0.5300 1.8360 0.5420 ;
        RECT 1.7860 0.5420 1.8360 0.9560 ;
        RECT 1.6470 0.4920 1.9110 0.5300 ;
        RECT 1.6470 0.9560 1.8360 1.0060 ;
        RECT 1.7510 0.3920 1.9110 0.4920 ;
        RECT 1.6470 0.1880 1.6970 0.4920 ;
        RECT 1.6470 1.0060 1.6970 1.4260 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN A5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0230 0.5410 1.1230 0.5490 ;
        RECT 1.0090 0.5490 1.1230 0.6010 ;
        RECT 1.0090 0.6010 1.1650 0.6750 ;
        RECT 1.1150 0.6750 1.1650 0.8080 ;
    END
    ANTENNAGATEAREA 0.0231 ;
  END A5
  OBS
    LAYER NWELL ;
      RECT -0.1350 0.6790 2.0920 1.7870 ;
    LAYER M1 ;
      RECT 1.3430 0.6310 1.6210 0.6810 ;
      RECT 1.5350 0.6810 1.6210 0.6990 ;
      RECT 1.5350 0.6130 1.6210 0.6310 ;
      RECT 1.3430 0.5330 1.3930 0.6310 ;
      RECT 1.3430 0.6810 1.3930 0.9030 ;
      RECT 1.1910 0.4830 1.3930 0.5330 ;
      RECT 1.0390 0.9030 1.3930 0.9530 ;
      RECT 1.1910 0.2110 1.2410 0.4830 ;
      RECT 1.3430 0.9530 1.3930 1.3800 ;
      RECT 1.0390 0.9530 1.0890 1.2130 ;
      RECT 0.5830 1.2130 1.0890 1.2630 ;
      RECT 0.5830 1.2630 0.6330 1.3930 ;
      RECT 0.5830 1.1060 0.6330 1.2130 ;
      RECT 0.2790 0.5980 0.9370 0.6480 ;
      RECT 0.8870 0.2080 0.9370 0.5980 ;
      RECT 0.5830 0.1810 0.6330 0.5980 ;
      RECT 0.2790 0.1780 0.3290 0.5980 ;
      RECT 1.3430 0.1480 1.3930 0.4320 ;
      RECT 0.7350 0.0980 1.3930 0.1480 ;
      RECT 1.0390 0.1480 1.0890 0.4310 ;
      RECT 0.7350 0.1480 0.7850 0.5010 ;
    LAYER PO ;
      RECT 1.2770 0.1010 1.3070 1.5670 ;
      RECT 1.5810 0.0690 1.6110 1.6080 ;
      RECT 1.1250 0.1010 1.1550 1.4690 ;
      RECT 1.4290 0.1010 1.4590 1.4690 ;
      RECT 0.3650 0.1010 0.3950 1.4690 ;
      RECT 1.8850 0.1010 1.9150 1.4690 ;
      RECT 0.0610 0.1010 0.0910 1.4690 ;
      RECT 1.7330 0.1010 1.7630 1.4690 ;
      RECT 0.9730 0.1010 1.0030 1.4690 ;
      RECT 0.8210 0.1010 0.8510 1.4690 ;
      RECT 0.6690 0.1010 0.6990 1.4690 ;
      RECT 0.5170 0.1010 0.5470 1.5670 ;
      RECT 0.2130 0.1010 0.2430 1.4690 ;
  END
END OA222X1_LVT

MACRO OA222X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.128 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.1280 0.0300 ;
        RECT 0.4310 0.0300 0.4810 0.5120 ;
        RECT 1.6470 0.0300 1.6970 0.3990 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7100 0.4210 0.8170 ;
        RECT 0.2490 0.7010 0.3590 0.7100 ;
    END
    ANTENNAGATEAREA 0.0231 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 1.4610 0.5730 1.5750 ;
        RECT 0.4260 1.4600 0.5730 1.4610 ;
    END
    ANTENNAGATEAREA 0.0231 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8110 0.7720 0.8610 1.0020 ;
        RECT 0.8110 1.0020 0.9680 1.1390 ;
    END
    ANTENNAGATEAREA 0.0231 ;
  END A3

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6590 0.7130 0.7090 0.8540 ;
        RECT 0.5530 0.8540 0.7090 0.9860 ;
    END
    ANTENNAGATEAREA 0.0231 ;
  END A4

  PIN A5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0230 0.5410 1.1230 0.5490 ;
        RECT 1.0090 0.5490 1.1230 0.6010 ;
        RECT 1.0090 0.6010 1.1650 0.6580 ;
        RECT 1.0230 0.6580 1.1650 0.6750 ;
        RECT 1.1150 0.6750 1.1650 0.8080 ;
    END
    ANTENNAGATEAREA 0.0231 ;
  END A5

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9380 0.5420 1.9880 0.9560 ;
        RECT 1.4950 0.5300 1.9880 0.5420 ;
        RECT 1.4950 0.9560 1.9880 1.0060 ;
        RECT 1.4950 0.4920 2.0630 0.5300 ;
        RECT 1.7990 1.0060 1.8490 1.4260 ;
        RECT 1.4950 1.0060 1.5450 1.4260 ;
        RECT 1.9030 0.3920 2.0630 0.4920 ;
        RECT 1.7990 0.1880 1.8490 0.4920 ;
        RECT 1.4950 0.1880 1.5450 0.4920 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END Y

  PIN A6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1600 1.1460 1.2800 1.2810 ;
        RECT 1.1710 1.2810 1.2210 1.4850 ;
        RECT 1.1710 1.4850 1.3390 1.5350 ;
    END
    ANTENNAGATEAREA 0.0231 ;
  END A6

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.1280 1.7020 ;
        RECT 0.8870 1.3350 0.9370 1.6420 ;
        RECT 1.0390 1.3330 1.0890 1.6420 ;
        RECT 0.2790 0.9580 0.3290 1.6420 ;
        RECT 1.6470 1.1330 1.6970 1.6420 ;
    END
  END VDD
  OBS
    LAYER NWELL ;
      RECT -0.1350 0.6790 2.2440 1.7870 ;
    LAYER M1 ;
      RECT 1.6870 0.6810 1.7730 0.6990 ;
      RECT 1.3430 0.6310 1.7730 0.6810 ;
      RECT 1.6870 0.6130 1.7730 0.6310 ;
      RECT 1.5260 0.6810 1.6120 0.6990 ;
      RECT 1.5260 0.6130 1.6120 0.6310 ;
      RECT 0.5830 1.2630 0.6330 1.3930 ;
      RECT 0.5830 1.1060 0.6330 1.2130 ;
      RECT 1.3430 0.6810 1.3930 0.9030 ;
      RECT 1.3430 0.5330 1.3930 0.6310 ;
      RECT 1.0390 0.9030 1.3930 0.9530 ;
      RECT 1.1910 0.4830 1.3930 0.5330 ;
      RECT 1.3430 0.9530 1.3930 1.3800 ;
      RECT 1.1910 0.2110 1.2410 0.4830 ;
      RECT 1.0390 0.9530 1.0890 1.2130 ;
      RECT 0.5830 1.2130 1.0890 1.2630 ;
      RECT 1.0390 0.1480 1.0890 0.4310 ;
      RECT 0.7350 0.0980 1.3930 0.1480 ;
      RECT 1.3430 0.1480 1.3930 0.4320 ;
      RECT 0.7350 0.1480 0.7850 0.5010 ;
      RECT 0.2790 0.5980 0.9370 0.6480 ;
      RECT 0.5830 0.1810 0.6330 0.5980 ;
      RECT 0.8870 0.2080 0.9370 0.5980 ;
      RECT 0.2790 0.1780 0.3290 0.5980 ;
    LAYER PO ;
      RECT 1.5810 0.0690 1.6110 1.6080 ;
      RECT 1.7330 0.0690 1.7630 1.6080 ;
      RECT 0.8210 0.1010 0.8510 1.4690 ;
      RECT 0.6690 0.1010 0.6990 1.4690 ;
      RECT 0.5170 0.1010 0.5470 1.5670 ;
      RECT 0.2130 0.1010 0.2430 1.4690 ;
      RECT 1.2770 0.1010 1.3070 1.5670 ;
      RECT 1.1250 0.1010 1.1550 1.4690 ;
      RECT 0.3650 0.1010 0.3950 1.4690 ;
      RECT 1.4290 0.1010 1.4590 1.4690 ;
      RECT 1.8850 0.1010 1.9150 1.4690 ;
      RECT 2.0370 0.1010 2.0670 1.4690 ;
      RECT 0.0610 0.1010 0.0910 1.4690 ;
      RECT 0.9730 0.1010 1.0030 1.4690 ;
  END
END OA222X2_LVT

MACRO OA22X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.52 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.5200 1.7020 ;
        RECT 0.8870 1.3350 0.9370 1.6420 ;
        RECT 0.2790 0.9580 0.3290 1.6420 ;
        RECT 1.0390 1.3330 1.0890 1.6420 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3300 0.5420 1.3800 0.9560 ;
        RECT 1.1910 0.5300 1.3800 0.5420 ;
        RECT 1.1910 0.9560 1.3800 1.0060 ;
        RECT 1.1910 0.4920 1.4550 0.5300 ;
        RECT 1.1910 1.0060 1.2410 1.4260 ;
        RECT 1.2950 0.3920 1.4550 0.4920 ;
        RECT 1.1910 0.1880 1.2410 0.4920 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6590 0.7230 0.7090 0.8540 ;
        RECT 0.5530 0.8540 0.7090 0.9860 ;
    END
    ANTENNAGATEAREA 0.0216 ;
  END A4

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8110 0.7150 0.8610 1.0020 ;
        RECT 0.8110 1.0020 0.9680 1.1390 ;
    END
    ANTENNAGATEAREA 0.0216 ;
  END A3

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 1.4610 0.5730 1.5750 ;
        RECT 0.4260 1.4600 0.5730 1.4610 ;
    END
    ANTENNAGATEAREA 0.0216 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7010 0.3590 0.7100 ;
        RECT 0.2490 0.7100 0.4210 0.8100 ;
        RECT 0.2710 0.8100 0.4210 0.8170 ;
    END
    ANTENNAGATEAREA 0.0216 ;
  END A1

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.5200 0.0300 ;
        RECT 0.4310 0.0300 0.4810 0.5120 ;
        RECT 1.0390 0.0300 1.0890 0.3990 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1350 0.6790 1.6360 1.7870 ;
    LAYER M1 ;
      RECT 1.0790 0.6630 1.1650 0.6990 ;
      RECT 0.7350 0.6130 1.1650 0.6630 ;
      RECT 1.0790 0.6990 1.1290 1.2260 ;
      RECT 0.5830 1.2260 1.1290 1.2760 ;
      RECT 0.7350 0.2120 0.7850 0.6130 ;
      RECT 0.5830 1.2760 0.6330 1.3930 ;
      RECT 0.5830 1.1060 0.6330 1.2260 ;
      RECT 0.5830 0.0950 0.9370 0.1450 ;
      RECT 0.5830 0.1450 0.6330 0.5980 ;
      RECT 0.8870 0.1450 0.9370 0.5040 ;
      RECT 0.2790 0.5980 0.6330 0.6480 ;
      RECT 0.2790 0.1780 0.3290 0.5980 ;
    LAYER PO ;
      RECT 0.0610 0.1010 0.0910 1.4690 ;
      RECT 0.5170 0.1010 0.5470 1.5670 ;
      RECT 0.2130 0.1010 0.2430 1.4690 ;
      RECT 0.9730 0.1010 1.0030 1.4690 ;
      RECT 0.8210 0.1010 0.8510 1.4690 ;
      RECT 0.6690 0.1010 0.6990 1.4690 ;
      RECT 1.1250 0.0690 1.1550 1.6080 ;
      RECT 0.3650 0.1010 0.3950 1.4690 ;
      RECT 1.2770 0.1010 1.3070 1.4690 ;
      RECT 1.4290 0.1010 1.4590 1.4690 ;
  END
END OA22X1_LVT

MACRO OA22X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.672 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.6720 1.7020 ;
        RECT 0.2790 0.9580 0.3290 1.6420 ;
        RECT 0.8870 1.3350 0.9370 1.6420 ;
        RECT 1.1910 1.4610 1.2410 1.6420 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0390 0.5300 1.5320 0.5420 ;
        RECT 1.4820 0.5420 1.5320 0.9560 ;
        RECT 1.0390 0.4920 1.6070 0.5300 ;
        RECT 1.3430 0.9560 1.5320 1.0060 ;
        RECT 1.4470 0.3920 1.6070 0.4920 ;
        RECT 1.3430 0.1880 1.3930 0.4920 ;
        RECT 1.0390 0.1880 1.0890 0.4920 ;
        RECT 1.3430 1.0060 1.3930 1.3390 ;
        RECT 1.0390 1.3390 1.3930 1.3890 ;
        RECT 1.0390 1.3890 1.0890 1.5580 ;
        RECT 1.3430 1.3890 1.3930 1.4260 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END Y

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6590 0.7230 0.7090 0.8540 ;
        RECT 0.5530 0.8540 0.7090 0.9860 ;
    END
    ANTENNAGATEAREA 0.0216 ;
  END A4

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8110 0.7150 0.8610 1.0020 ;
        RECT 0.8110 1.0020 0.9680 1.1390 ;
    END
    ANTENNAGATEAREA 0.0216 ;
  END A3

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 1.4610 0.5730 1.5750 ;
        RECT 0.4260 1.4600 0.5730 1.4610 ;
    END
    ANTENNAGATEAREA 0.0216 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7010 0.3590 0.7100 ;
        RECT 0.2490 0.7100 0.4210 0.8170 ;
    END
    ANTENNAGATEAREA 0.0216 ;
  END A1

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.6720 0.0300 ;
        RECT 0.4310 0.0300 0.4810 0.5120 ;
        RECT 1.1910 0.0300 1.2410 0.3990 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1350 0.6790 1.7880 1.7870 ;
    LAYER M1 ;
      RECT 1.2310 0.6810 1.3170 0.6990 ;
      RECT 1.0700 0.6630 1.3170 0.6810 ;
      RECT 0.7350 0.6310 1.3170 0.6630 ;
      RECT 1.2310 0.6130 1.3170 0.6310 ;
      RECT 1.0700 0.6810 1.1560 0.6990 ;
      RECT 0.7350 0.6130 1.1560 0.6310 ;
      RECT 0.7350 0.2120 0.7850 0.6130 ;
      RECT 1.0790 0.6990 1.1290 1.2260 ;
      RECT 0.5830 1.2260 1.1290 1.2760 ;
      RECT 0.5830 1.2760 0.6330 1.3930 ;
      RECT 0.5830 1.1060 0.6330 1.2260 ;
      RECT 0.5830 0.0950 0.9370 0.1450 ;
      RECT 0.8870 0.1450 0.9370 0.5040 ;
      RECT 0.5830 0.1450 0.6330 0.5980 ;
      RECT 0.2790 0.5980 0.6330 0.6480 ;
      RECT 0.2790 0.1780 0.3290 0.5980 ;
    LAYER PO ;
      RECT 1.4290 0.1010 1.4590 1.4690 ;
      RECT 0.8210 0.1010 0.8510 1.4690 ;
      RECT 0.6690 0.1010 0.6990 1.4690 ;
      RECT 1.1250 0.0690 1.1550 1.6080 ;
      RECT 0.3650 0.1010 0.3950 1.4690 ;
      RECT 1.5810 0.1010 1.6110 1.4690 ;
      RECT 0.5170 0.1010 0.5470 1.5670 ;
      RECT 1.2770 0.0690 1.3070 1.6080 ;
      RECT 0.9730 0.1010 1.0030 1.4690 ;
      RECT 0.0610 0.1010 0.0910 1.4690 ;
      RECT 0.2130 0.1010 0.2430 1.4690 ;
  END
END OA22X2_LVT

MACRO OAI21X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.824 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.8240 1.7020 ;
        RECT 0.2790 0.9580 0.3290 1.6420 ;
        RECT 1.0390 1.4140 1.0890 1.6420 ;
        RECT 0.8870 1.2430 0.9370 1.6420 ;
        RECT 1.3430 1.1330 1.3930 1.6420 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6340 0.5420 1.6840 0.9560 ;
        RECT 1.4950 0.5300 1.6840 0.5420 ;
        RECT 1.4950 0.9560 1.6840 1.0060 ;
        RECT 1.4950 0.4920 1.7430 0.5300 ;
        RECT 1.4950 1.0060 1.5450 1.4260 ;
        RECT 1.6070 0.3920 1.7430 0.4920 ;
        RECT 1.4950 0.1880 1.5450 0.4920 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 0.8530 0.8610 0.9620 ;
        RECT 0.7120 0.9620 0.8610 0.9860 ;
        RECT 0.8110 0.8070 0.8610 0.8530 ;
    END
    ANTENNAGATEAREA 0.0138 ;
  END A3

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4000 1.4610 0.5730 1.5750 ;
        RECT 0.4260 1.4600 0.5730 1.4610 ;
    END
    ANTENNAGATEAREA 0.0246 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7010 0.3590 0.7170 ;
        RECT 0.2490 0.7170 0.4210 0.8150 ;
        RECT 0.2710 0.8150 0.4210 0.8170 ;
    END
    ANTENNAGATEAREA 0.0246 ;
  END A1

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.8240 0.0300 ;
        RECT 0.4310 0.0300 0.4810 0.5120 ;
        RECT 1.0390 0.0300 1.0890 0.2340 ;
        RECT 1.3430 0.0300 1.3930 0.3990 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1140 0.6790 1.9390 1.7870 ;
    LAYER M1 ;
      RECT 1.0790 0.7850 1.1650 0.8030 ;
      RECT 0.9130 0.7550 1.1650 0.7850 ;
      RECT 0.8870 0.7350 1.1650 0.7550 ;
      RECT 1.0790 0.7170 1.1650 0.7350 ;
      RECT 0.7350 1.1800 0.7850 1.3930 ;
      RECT 0.9130 0.7850 0.9630 1.1300 ;
      RECT 0.8870 0.7050 0.9630 0.7350 ;
      RECT 0.5830 1.1300 0.9630 1.1800 ;
      RECT 0.8870 0.1810 0.9370 0.7050 ;
      RECT 0.5830 1.1800 0.6330 1.3930 ;
      RECT 0.5830 1.1060 0.6330 1.1300 ;
      RECT 1.2310 0.6310 1.4800 0.6810 ;
      RECT 1.3830 0.6810 1.4690 0.6990 ;
      RECT 1.3830 0.6130 1.4690 0.6310 ;
      RECT 1.2310 0.6810 1.2810 0.9560 ;
      RECT 1.2310 0.5420 1.2810 0.6310 ;
      RECT 1.1910 0.9560 1.2810 1.0060 ;
      RECT 1.1910 0.4920 1.2810 0.5420 ;
      RECT 1.1910 1.0060 1.2410 1.5550 ;
      RECT 1.1910 0.0880 1.2410 0.4920 ;
      RECT 0.2790 0.5980 0.6330 0.6480 ;
      RECT 0.5830 0.4620 0.6330 0.5980 ;
      RECT 0.5830 0.4120 0.7850 0.4620 ;
      RECT 0.7350 0.1810 0.7850 0.4120 ;
      RECT 0.5830 0.1810 0.6330 0.4120 ;
      RECT 0.2790 0.1780 0.3290 0.5980 ;
    LAYER PO ;
      RECT 0.9730 0.1010 1.0030 1.4690 ;
      RECT 1.1250 0.0540 1.1550 1.6080 ;
      RECT 0.3650 0.1010 0.3950 1.4690 ;
      RECT 0.8210 0.1010 0.8510 1.4690 ;
      RECT 1.5810 0.1010 1.6110 1.4690 ;
      RECT 1.7330 0.1010 1.7630 1.4690 ;
      RECT 0.0610 0.1010 0.0910 1.4690 ;
      RECT 1.2770 0.1010 1.3070 1.4690 ;
      RECT 1.4290 0.0690 1.4590 1.6080 ;
      RECT 0.5170 0.1010 0.5470 1.5670 ;
      RECT 0.2130 0.1010 0.2430 1.4690 ;
      RECT 0.6690 0.1010 0.6990 1.4690 ;
  END
END OAI21X1_LVT

MACRO OAI21X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.976 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.9760 1.7020 ;
        RECT 0.2790 0.9580 0.3290 1.6420 ;
        RECT 1.0390 1.4140 1.0890 1.6420 ;
        RECT 0.8870 1.2430 0.9370 1.6420 ;
        RECT 1.4950 1.1330 1.5450 1.6420 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3430 0.5300 1.8360 0.5420 ;
        RECT 1.7860 0.5420 1.8360 0.9560 ;
        RECT 1.3430 0.4920 1.8950 0.5300 ;
        RECT 1.3430 0.9560 1.8360 1.0060 ;
        RECT 1.7590 0.3920 1.8950 0.4920 ;
        RECT 1.6470 0.1880 1.6970 0.4920 ;
        RECT 1.3430 0.1880 1.3930 0.4920 ;
        RECT 1.6470 1.0060 1.6970 1.4260 ;
        RECT 1.3430 1.0060 1.3930 1.4260 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END Y

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 0.8530 0.8610 0.9670 ;
        RECT 0.7120 0.9670 0.8610 0.9860 ;
        RECT 0.8110 0.8070 0.8610 0.8530 ;
    END
    ANTENNAGATEAREA 0.0156 ;
  END A3

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4000 1.4610 0.5730 1.5750 ;
        RECT 0.4260 1.4600 0.5730 1.4610 ;
    END
    ANTENNAGATEAREA 0.0258 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7010 0.3590 0.7170 ;
        RECT 0.2490 0.7170 0.4210 0.8150 ;
        RECT 0.2710 0.8150 0.4210 0.8170 ;
    END
    ANTENNAGATEAREA 0.0258 ;
  END A1

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.9760 0.0300 ;
        RECT 0.4310 0.0300 0.4810 0.5120 ;
        RECT 1.0390 0.0300 1.0890 0.2340 ;
        RECT 1.4950 0.0300 1.5450 0.3990 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 2.0910 1.7870 ;
    LAYER M1 ;
      RECT 1.0790 0.7850 1.1650 0.8030 ;
      RECT 0.9130 0.7550 1.1650 0.7850 ;
      RECT 0.8870 0.7350 1.1650 0.7550 ;
      RECT 1.0790 0.7170 1.1650 0.7350 ;
      RECT 0.7350 1.1800 0.7850 1.3930 ;
      RECT 0.7350 1.1060 0.7850 1.1300 ;
      RECT 0.9130 0.7850 0.9630 1.1300 ;
      RECT 0.8870 0.7050 0.9630 0.7350 ;
      RECT 0.5830 1.1300 0.9630 1.1800 ;
      RECT 0.8870 0.1810 0.9370 0.7050 ;
      RECT 0.5830 1.1800 0.6330 1.3930 ;
      RECT 0.5830 1.1060 0.6330 1.1300 ;
      RECT 1.5350 0.6810 1.6210 0.6990 ;
      RECT 1.2310 0.6310 1.6210 0.6810 ;
      RECT 1.5350 0.6130 1.6210 0.6310 ;
      RECT 1.3740 0.6810 1.4600 0.6990 ;
      RECT 1.3740 0.6130 1.4600 0.6310 ;
      RECT 1.2310 0.6810 1.2810 0.9560 ;
      RECT 1.2310 0.5420 1.2810 0.6310 ;
      RECT 1.1910 0.9560 1.2810 1.0060 ;
      RECT 1.1910 0.4920 1.2810 0.5420 ;
      RECT 1.1910 1.0060 1.2410 1.5550 ;
      RECT 1.1910 0.0960 1.2410 0.4920 ;
      RECT 0.2790 0.5980 0.6330 0.6480 ;
      RECT 0.5830 0.4620 0.6330 0.5980 ;
      RECT 0.5830 0.4120 0.7850 0.4620 ;
      RECT 0.7350 0.1810 0.7850 0.4120 ;
      RECT 0.5830 0.1810 0.6330 0.4120 ;
      RECT 0.2790 0.1780 0.3290 0.5980 ;
    LAYER PO ;
      RECT 0.9730 0.1010 1.0030 1.4690 ;
      RECT 1.1250 0.0540 1.1550 1.6080 ;
      RECT 1.4290 0.0690 1.4590 1.6080 ;
      RECT 0.3650 0.1010 0.3950 1.4690 ;
      RECT 0.8210 0.1010 0.8510 1.4690 ;
      RECT 1.7330 0.1010 1.7630 1.4690 ;
      RECT 1.8850 0.1010 1.9150 1.4690 ;
      RECT 0.0610 0.1010 0.0910 1.4690 ;
      RECT 1.2770 0.1010 1.3070 1.4690 ;
      RECT 1.5810 0.0690 1.6110 1.6080 ;
      RECT 0.5170 0.1010 0.5470 1.5670 ;
      RECT 0.2130 0.1010 0.2430 1.4690 ;
      RECT 0.6690 0.1010 0.6990 1.4690 ;
  END
END OAI21X2_LVT

MACRO OAI221X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.128 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7990 0.5300 1.9880 0.5420 ;
        RECT 1.9380 0.5420 1.9880 0.9560 ;
        RECT 1.7990 0.4920 2.0630 0.5300 ;
        RECT 1.7990 0.9560 1.9880 1.0060 ;
        RECT 1.9030 0.3920 2.0630 0.4920 ;
        RECT 1.7990 0.1880 1.8490 0.4920 ;
        RECT 1.7990 1.0060 1.8490 1.4260 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN A5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0230 0.5410 1.1230 0.5490 ;
        RECT 1.0090 0.5490 1.1230 0.6010 ;
        RECT 1.0090 0.6010 1.1650 0.6630 ;
        RECT 1.0230 0.6630 1.1650 0.6750 ;
        RECT 1.1150 0.6750 1.1650 0.8080 ;
    END
    ANTENNAGATEAREA 0.0162 ;
  END A5

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7010 0.3590 0.7100 ;
        RECT 0.2490 0.7100 0.4210 0.8150 ;
        RECT 0.2710 0.8150 0.4210 0.8170 ;
    END
    ANTENNAGATEAREA 0.0222 ;
  END A1

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.1280 0.0300 ;
        RECT 1.6470 0.0300 1.6970 0.3990 ;
        RECT 1.3430 0.0300 1.3930 0.5320 ;
        RECT 0.4310 0.0300 0.4810 0.5120 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.1280 1.7020 ;
        RECT 1.0390 1.3330 1.0890 1.6420 ;
        RECT 1.3430 1.2340 1.3930 1.6420 ;
        RECT 1.6470 1.1330 1.6970 1.6420 ;
        RECT 0.2790 0.9580 0.3290 1.6420 ;
        RECT 0.8870 1.3350 0.9370 1.6420 ;
    END
  END VDD

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 0.8540 0.7090 0.9670 ;
        RECT 0.5600 0.9670 0.7090 0.9860 ;
        RECT 0.6590 0.7130 0.7090 0.8540 ;
    END
    ANTENNAGATEAREA 0.0222 ;
  END A4

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8110 0.8420 0.8610 1.0020 ;
        RECT 0.8110 1.0020 0.9680 1.1390 ;
    END
    ANTENNAGATEAREA 0.0222 ;
  END A3

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 1.4650 0.5110 1.4780 ;
        RECT 0.4010 1.4780 0.5730 1.5280 ;
        RECT 0.4010 1.5280 0.5110 1.5750 ;
    END
    ANTENNAGATEAREA 0.0222 ;
  END A2
  OBS
    LAYER NWELL ;
      RECT -0.1140 0.6790 2.2440 1.7870 ;
    LAYER M1 ;
      RECT 1.6870 0.6810 1.7730 0.6990 ;
      RECT 1.5350 0.6310 1.7730 0.6810 ;
      RECT 1.6870 0.6130 1.7730 0.6310 ;
      RECT 1.5350 0.6810 1.5850 0.9560 ;
      RECT 1.5350 0.5420 1.5850 0.6310 ;
      RECT 1.4950 0.9560 1.5850 1.0060 ;
      RECT 1.4950 0.4920 1.5850 0.5420 ;
      RECT 1.4950 1.0060 1.5450 1.4260 ;
      RECT 1.4950 0.1880 1.5450 0.4920 ;
      RECT 1.0390 0.9030 1.4320 0.9530 ;
      RECT 1.3820 0.8030 1.4320 0.9030 ;
      RECT 1.3820 0.7170 1.4690 0.8030 ;
      RECT 1.1910 0.9530 1.2410 1.4270 ;
      RECT 1.2270 0.5330 1.2770 0.9030 ;
      RECT 1.0390 0.9530 1.0890 1.2130 ;
      RECT 1.1910 0.4830 1.2770 0.5330 ;
      RECT 0.5830 1.2130 1.0890 1.2630 ;
      RECT 1.1910 0.2110 1.2410 0.4830 ;
      RECT 0.5830 1.2630 0.6330 1.3930 ;
      RECT 0.5830 1.1060 0.6330 1.2130 ;
      RECT 0.2790 0.5980 0.9370 0.6480 ;
      RECT 0.8870 0.2080 0.9370 0.5980 ;
      RECT 0.5830 0.1810 0.6330 0.5980 ;
      RECT 0.2790 0.1780 0.3290 0.5980 ;
      RECT 0.7350 0.0980 1.0890 0.1480 ;
      RECT 1.0390 0.1480 1.0890 0.4310 ;
      RECT 0.7350 0.1480 0.7850 0.5010 ;
    LAYER PO ;
      RECT 0.9730 0.1010 1.0030 1.4690 ;
      RECT 0.0610 0.1010 0.0910 1.4690 ;
      RECT 2.0370 0.1010 2.0670 1.4690 ;
      RECT 1.8850 0.1010 1.9150 1.4690 ;
      RECT 1.2770 0.1010 1.3070 1.4690 ;
      RECT 0.3650 0.1010 0.3950 1.4690 ;
      RECT 1.5810 0.1010 1.6110 1.4690 ;
      RECT 1.1250 0.1010 1.1550 1.4690 ;
      RECT 1.7330 0.0690 1.7630 1.6080 ;
      RECT 0.2130 0.1010 0.2430 1.4690 ;
      RECT 0.5170 0.1010 0.5470 1.5670 ;
      RECT 1.4290 0.0540 1.4590 1.6080 ;
      RECT 0.6690 0.1010 0.6990 1.4690 ;
      RECT 0.8210 0.1010 0.8510 1.4690 ;
  END
END OAI221X1_LVT

MACRO OAI221X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.28 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.2800 1.7020 ;
        RECT 0.2790 0.9580 0.3290 1.6420 ;
        RECT 1.7990 1.1330 1.8490 1.6420 ;
        RECT 1.3430 1.2340 1.3930 1.6420 ;
        RECT 0.8870 1.3350 0.9370 1.6420 ;
        RECT 1.0390 1.3330 1.0890 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.2800 0.0300 ;
        RECT 0.4310 0.0300 0.4810 0.5120 ;
        RECT 1.7990 0.0300 1.8490 0.3990 ;
        RECT 1.3430 0.0300 1.3930 0.5320 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7010 0.3590 0.7100 ;
        RECT 0.2490 0.7100 0.4210 0.8150 ;
        RECT 0.2710 0.8150 0.4210 0.8170 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END A1

  PIN A5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0230 0.5410 1.1230 0.5490 ;
        RECT 1.0090 0.5490 1.1230 0.6010 ;
        RECT 1.0090 0.6010 1.1650 0.6630 ;
        RECT 1.0230 0.6630 1.1650 0.6750 ;
        RECT 1.1150 0.6750 1.1650 0.8080 ;
    END
    ANTENNAGATEAREA 0.0162 ;
  END A5

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6470 0.5300 2.1400 0.5420 ;
        RECT 2.0900 0.5420 2.1400 0.9560 ;
        RECT 1.6470 0.4920 2.2150 0.5300 ;
        RECT 1.6470 0.9560 2.1400 1.0060 ;
        RECT 2.0550 0.3920 2.2150 0.4920 ;
        RECT 1.9510 0.1880 2.0010 0.4920 ;
        RECT 1.6470 0.1880 1.6970 0.4920 ;
        RECT 1.9510 1.0060 2.0010 1.4260 ;
        RECT 1.6470 1.0060 1.6970 1.4260 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END Y

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 1.4610 0.5730 1.5750 ;
        RECT 0.4260 1.4600 0.5730 1.4610 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8110 0.8420 0.8610 1.0020 ;
        RECT 0.8110 1.0020 0.9680 1.1390 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END A3

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 0.8540 0.7090 0.9670 ;
        RECT 0.5600 0.9670 0.7090 0.9860 ;
        RECT 0.6590 0.7130 0.7090 0.8540 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END A4
  OBS
    LAYER NWELL ;
      RECT -0.1140 0.6790 2.3960 1.7870 ;
    LAYER M1 ;
      RECT 1.8390 0.6810 1.9250 0.6990 ;
      RECT 1.5350 0.6310 1.9250 0.6810 ;
      RECT 1.8390 0.6130 1.9250 0.6310 ;
      RECT 1.5350 0.6810 1.5850 0.9560 ;
      RECT 1.5350 0.5420 1.5850 0.6310 ;
      RECT 1.4950 0.9560 1.5850 1.0060 ;
      RECT 1.4950 0.4920 1.5850 0.5420 ;
      RECT 1.4950 1.0060 1.5450 1.4260 ;
      RECT 1.4950 0.1880 1.5450 0.4920 ;
      RECT 1.6870 0.6810 1.7730 0.6990 ;
      RECT 1.6870 0.6130 1.7730 0.6310 ;
      RECT 1.0390 0.9030 1.4320 0.9530 ;
      RECT 1.3820 0.8030 1.4320 0.9030 ;
      RECT 1.3820 0.7170 1.4690 0.8030 ;
      RECT 1.1910 0.9530 1.2410 1.4270 ;
      RECT 1.2270 0.5330 1.2770 0.9030 ;
      RECT 1.0390 0.9530 1.0890 1.2130 ;
      RECT 1.1910 0.4830 1.2770 0.5330 ;
      RECT 0.5830 1.2130 1.0890 1.2630 ;
      RECT 1.1910 0.2110 1.2410 0.4830 ;
      RECT 0.5830 1.2630 0.6330 1.3930 ;
      RECT 0.5830 1.1060 0.6330 1.2130 ;
      RECT 0.2790 0.5980 0.9370 0.6480 ;
      RECT 0.5830 0.1810 0.6330 0.5980 ;
      RECT 0.8870 0.2080 0.9370 0.5980 ;
      RECT 0.2790 0.1780 0.3290 0.5980 ;
      RECT 0.7350 0.0980 1.0890 0.1480 ;
      RECT 1.0390 0.1480 1.0890 0.4310 ;
      RECT 0.7350 0.1480 0.7850 0.5010 ;
    LAYER PO ;
      RECT 0.6690 0.1010 0.6990 1.4690 ;
      RECT 0.3650 0.1010 0.3950 1.4690 ;
      RECT 1.2770 0.1010 1.3070 1.4690 ;
      RECT 0.9730 0.1010 1.0030 1.4690 ;
      RECT 0.0610 0.1010 0.0910 1.4690 ;
      RECT 0.2130 0.1010 0.2430 1.4690 ;
      RECT 2.0370 0.1010 2.0670 1.4690 ;
      RECT 0.8210 0.1010 0.8510 1.4690 ;
      RECT 1.5810 0.1010 1.6110 1.4690 ;
      RECT 1.1250 0.1010 1.1550 1.4690 ;
      RECT 2.1890 0.1010 2.2190 1.4690 ;
      RECT 0.5170 0.1010 0.5470 1.5670 ;
      RECT 1.8850 0.0690 1.9150 1.6080 ;
      RECT 1.4290 0.0540 1.4590 1.6080 ;
      RECT 1.7330 0.0690 1.7630 1.6080 ;
  END
END OAI221X2_LVT

MACRO OAI222X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.28 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.2800 1.7020 ;
        RECT 0.2790 0.9580 0.3290 1.6420 ;
        RECT 1.0390 1.3330 1.0890 1.6420 ;
        RECT 0.8870 1.3350 0.9370 1.6420 ;
        RECT 1.4950 1.2340 1.5450 1.6420 ;
        RECT 1.7990 1.1330 1.8490 1.6420 ;
    END
  END VDD

  PIN A6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1600 1.1460 1.2800 1.2810 ;
        RECT 1.1710 1.2810 1.2210 1.4850 ;
        RECT 1.1710 1.4850 1.3390 1.5350 ;
    END
    ANTENNAGATEAREA 0.0225 ;
  END A6

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9510 0.5300 2.1400 0.5420 ;
        RECT 2.0900 0.5420 2.1400 0.9560 ;
        RECT 1.9510 0.4920 2.2150 0.5300 ;
        RECT 1.9510 0.9560 2.1400 1.0060 ;
        RECT 2.0550 0.3920 2.2150 0.4920 ;
        RECT 1.9510 0.1880 2.0010 0.4920 ;
        RECT 1.9510 1.0060 2.0010 1.4260 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN A5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0230 0.5410 1.1230 0.5490 ;
        RECT 1.0090 0.5490 1.1230 0.6010 ;
        RECT 1.0090 0.6010 1.1650 0.6630 ;
        RECT 1.0230 0.6630 1.1650 0.6750 ;
        RECT 1.1150 0.6750 1.1650 0.8080 ;
    END
    ANTENNAGATEAREA 0.0225 ;
  END A5

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 0.8540 0.7090 0.9860 ;
        RECT 0.6590 0.7130 0.7090 0.8540 ;
    END
    ANTENNAGATEAREA 0.0225 ;
  END A4

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8110 0.8420 0.8610 1.0020 ;
        RECT 0.8110 1.0020 0.9680 1.1390 ;
    END
    ANTENNAGATEAREA 0.0225 ;
  END A3

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 1.4610 0.5730 1.5750 ;
        RECT 0.4260 1.4600 0.5730 1.4610 ;
    END
    ANTENNAGATEAREA 0.0225 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7100 0.4210 0.8150 ;
        RECT 0.2490 0.7010 0.3590 0.7100 ;
        RECT 0.2710 0.8150 0.4210 0.8170 ;
    END
    ANTENNAGATEAREA 0.0225 ;
  END A1

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.2800 0.0300 ;
        RECT 0.4310 0.0300 0.4810 0.5120 ;
        RECT 1.4950 0.0300 1.5450 0.5320 ;
        RECT 1.7990 0.0300 1.8490 0.3990 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1370 0.6790 2.3940 1.7870 ;
    LAYER M1 ;
      RECT 1.8390 0.6810 1.9250 0.6990 ;
      RECT 1.6870 0.6310 1.9250 0.6810 ;
      RECT 1.8390 0.6130 1.9250 0.6310 ;
      RECT 1.6870 0.6810 1.7370 0.9560 ;
      RECT 1.6870 0.5420 1.7370 0.6310 ;
      RECT 1.6470 0.9560 1.7370 1.0060 ;
      RECT 1.6470 0.4920 1.7370 0.5420 ;
      RECT 1.6470 1.0060 1.6970 1.4260 ;
      RECT 1.6470 0.1880 1.6970 0.4920 ;
      RECT 1.5350 0.7170 1.6210 0.8030 ;
      RECT 1.5360 0.8030 1.5860 0.9030 ;
      RECT 1.0390 0.9030 1.5860 0.9530 ;
      RECT 1.3430 0.5330 1.3930 0.9030 ;
      RECT 1.3430 0.9530 1.3930 1.3800 ;
      RECT 1.1910 0.4830 1.3930 0.5330 ;
      RECT 1.1910 0.2110 1.2410 0.4830 ;
      RECT 1.0390 0.9530 1.0890 1.2130 ;
      RECT 0.5830 1.2130 1.0890 1.2630 ;
      RECT 0.5830 1.2630 0.6330 1.3930 ;
      RECT 0.5830 1.1060 0.6330 1.2130 ;
      RECT 0.2790 0.5980 0.9370 0.6480 ;
      RECT 0.8870 0.2080 0.9370 0.5980 ;
      RECT 0.5830 0.1810 0.6330 0.5980 ;
      RECT 0.2790 0.1780 0.3290 0.5980 ;
      RECT 1.0390 0.1480 1.0890 0.4310 ;
      RECT 0.7350 0.0980 1.3930 0.1480 ;
      RECT 1.3430 0.1480 1.3930 0.4320 ;
      RECT 0.7350 0.1480 0.7850 0.5010 ;
    LAYER PO ;
      RECT 0.6690 0.1010 0.6990 1.4690 ;
      RECT 0.8210 0.1010 0.8510 1.4690 ;
      RECT 2.0370 0.1010 2.0670 1.4690 ;
      RECT 0.2130 0.1010 0.2430 1.4690 ;
      RECT 0.0610 0.1010 0.0910 1.4690 ;
      RECT 0.9730 0.1010 1.0030 1.4690 ;
      RECT 1.4290 0.1010 1.4590 1.4690 ;
      RECT 0.3650 0.1010 0.3950 1.4690 ;
      RECT 1.7330 0.1010 1.7630 1.4690 ;
      RECT 1.1250 0.1010 1.1550 1.4690 ;
      RECT 2.1890 0.1010 2.2190 1.4690 ;
      RECT 0.5170 0.1010 0.5470 1.5670 ;
      RECT 1.2770 0.1010 1.3070 1.5670 ;
      RECT 1.8850 0.0690 1.9150 1.6080 ;
      RECT 1.5810 0.0540 1.6110 1.6080 ;
  END
END OAI222X1_LVT

MACRO OAI222X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.432 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.4320 1.7020 ;
        RECT 1.9510 1.1330 2.0010 1.6420 ;
        RECT 1.4950 1.2340 1.5450 1.6420 ;
        RECT 1.0390 1.3330 1.0890 1.6420 ;
        RECT 0.2790 0.9580 0.3290 1.6420 ;
        RECT 0.8870 1.3350 0.9370 1.6420 ;
    END
  END VDD

  PIN A6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1600 1.1570 1.2800 1.2710 ;
        RECT 1.1710 1.2710 1.2800 1.2810 ;
        RECT 1.1710 1.1460 1.2800 1.1570 ;
        RECT 1.1710 1.2810 1.2210 1.4850 ;
        RECT 1.1710 1.4850 1.3390 1.5350 ;
    END
    ANTENNAGATEAREA 0.0255 ;
  END A6

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7990 0.5300 2.2920 0.5420 ;
        RECT 2.2420 0.5420 2.2920 0.9560 ;
        RECT 1.7990 0.4920 2.3670 0.5300 ;
        RECT 1.7990 0.9560 2.2920 1.0060 ;
        RECT 2.2070 0.3920 2.3670 0.4920 ;
        RECT 2.1030 0.1880 2.1530 0.4920 ;
        RECT 1.7990 0.1880 1.8490 0.4920 ;
        RECT 2.1030 1.0060 2.1530 1.4260 ;
        RECT 1.7990 1.0060 1.8490 1.4260 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END Y

  PIN A5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0230 0.5410 1.1230 0.5490 ;
        RECT 1.0090 0.5490 1.1230 0.6010 ;
        RECT 1.0090 0.6010 1.1650 0.6630 ;
        RECT 1.0230 0.6630 1.1650 0.6750 ;
        RECT 1.1150 0.6750 1.1650 0.8080 ;
    END
    ANTENNAGATEAREA 0.0255 ;
  END A5

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5600 0.9630 0.7090 0.9860 ;
        RECT 0.5530 0.8540 0.7090 0.9630 ;
        RECT 0.6590 0.7130 0.7090 0.8540 ;
    END
    ANTENNAGATEAREA 0.0255 ;
  END A4

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8110 0.7720 0.8610 1.0020 ;
        RECT 0.8110 1.0020 0.9680 1.1390 ;
    END
    ANTENNAGATEAREA 0.0255 ;
  END A3

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 1.4610 0.5730 1.5750 ;
        RECT 0.4260 1.4600 0.5730 1.4610 ;
    END
    ANTENNAGATEAREA 0.0255 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7010 0.3590 0.7100 ;
        RECT 0.2490 0.7100 0.4210 0.8170 ;
    END
    ANTENNAGATEAREA 0.0255 ;
  END A1

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.4320 0.0300 ;
        RECT 1.9510 0.0300 2.0010 0.3990 ;
        RECT 1.4950 0.0300 1.5450 0.4040 ;
        RECT 0.4310 0.0300 0.4810 0.5120 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1110 0.6790 2.5480 1.7870 ;
    LAYER M1 ;
      RECT 1.9910 0.6810 2.0770 0.6990 ;
      RECT 1.6870 0.6310 2.0770 0.6810 ;
      RECT 1.9910 0.6130 2.0770 0.6310 ;
      RECT 1.8300 0.6810 1.9160 0.6990 ;
      RECT 1.8300 0.6130 1.9160 0.6310 ;
      RECT 1.6870 0.6810 1.7370 0.9560 ;
      RECT 1.6870 0.5420 1.7370 0.6310 ;
      RECT 1.6470 0.9560 1.7370 1.0060 ;
      RECT 1.6470 0.4920 1.7370 0.5420 ;
      RECT 1.6470 1.0060 1.6970 1.4260 ;
      RECT 1.6470 0.1880 1.6970 0.4920 ;
      RECT 1.5350 0.6640 1.6210 0.7500 ;
      RECT 1.5360 0.7500 1.5860 0.9030 ;
      RECT 1.0390 0.9030 1.5860 0.9530 ;
      RECT 1.3430 0.9530 1.3930 1.3800 ;
      RECT 1.3430 0.5330 1.3930 0.9030 ;
      RECT 1.1910 0.4830 1.3930 0.5330 ;
      RECT 1.1910 0.2110 1.2410 0.4830 ;
      RECT 1.0390 0.9530 1.0890 1.2130 ;
      RECT 0.5830 1.2130 1.0890 1.2630 ;
      RECT 0.5830 1.2630 0.6330 1.3930 ;
      RECT 0.5830 1.1060 0.6330 1.2130 ;
      RECT 1.0390 0.1480 1.0890 0.4310 ;
      RECT 0.7350 0.0980 1.3930 0.1480 ;
      RECT 1.3430 0.1480 1.3930 0.4320 ;
      RECT 0.7350 0.1480 0.7850 0.5010 ;
      RECT 0.2790 0.5980 0.9370 0.6480 ;
      RECT 0.8870 0.2080 0.9370 0.5980 ;
      RECT 0.5830 0.1810 0.6330 0.5980 ;
      RECT 0.2790 0.1780 0.3290 0.5980 ;
    LAYER PO ;
      RECT 1.8850 0.0690 1.9150 1.6080 ;
      RECT 0.6690 0.1010 0.6990 1.4690 ;
      RECT 0.8210 0.1010 0.8510 1.4690 ;
      RECT 2.3410 0.1010 2.3710 1.4690 ;
      RECT 1.5810 0.0540 1.6110 1.6080 ;
      RECT 0.5170 0.1010 0.5470 1.5670 ;
      RECT 0.2130 0.1010 0.2430 1.4690 ;
      RECT 2.0370 0.0690 2.0670 1.6080 ;
      RECT 1.1250 0.1010 1.1550 1.4690 ;
      RECT 1.7330 0.1010 1.7630 1.4690 ;
      RECT 0.3650 0.1010 0.3950 1.4690 ;
      RECT 1.4290 0.1010 1.4590 1.4690 ;
      RECT 2.1890 0.1010 2.2190 1.4690 ;
      RECT 0.0610 0.1010 0.0910 1.4690 ;
      RECT 1.2770 0.1010 1.3070 1.5670 ;
      RECT 0.9730 0.1010 1.0030 1.4690 ;
  END
END OAI222X2_LVT

MACRO OAI22X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.824 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.8240 1.7020 ;
        RECT 0.8870 1.3350 0.9370 1.6420 ;
        RECT 0.2790 0.9580 0.3290 1.6420 ;
        RECT 1.3430 1.1330 1.3930 1.6420 ;
        RECT 1.0390 1.3630 1.0890 1.6420 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6340 0.5420 1.6840 0.9560 ;
        RECT 1.4950 0.5300 1.6840 0.5420 ;
        RECT 1.4950 0.9560 1.6840 1.0060 ;
        RECT 1.4950 0.4920 1.7590 0.5300 ;
        RECT 1.4950 1.0060 1.5450 1.4260 ;
        RECT 1.5990 0.3920 1.7590 0.4920 ;
        RECT 1.4950 0.1880 1.5450 0.4920 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 0.8540 0.7090 0.9670 ;
        RECT 0.5600 0.9670 0.7090 0.9860 ;
        RECT 0.6590 0.7230 0.7090 0.8540 ;
    END
    ANTENNAGATEAREA 0.0276 ;
  END A4

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8110 0.7150 0.8610 1.0020 ;
        RECT 0.8110 1.0020 0.9680 1.1390 ;
    END
    ANTENNAGATEAREA 0.0276 ;
  END A3

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 1.4610 0.5730 1.5710 ;
        RECT 0.4010 1.5710 0.5110 1.5750 ;
        RECT 0.4260 1.4600 0.5730 1.4610 ;
    END
    ANTENNAGATEAREA 0.0276 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7010 0.3590 0.7100 ;
        RECT 0.2490 0.7100 0.4210 0.8150 ;
        RECT 0.2710 0.8150 0.4210 0.8170 ;
    END
    ANTENNAGATEAREA 0.0276 ;
  END A1

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.8240 0.0300 ;
        RECT 0.4310 0.0300 0.4810 0.5120 ;
        RECT 1.0390 0.0300 1.0890 0.4040 ;
        RECT 1.3430 0.0300 1.3930 0.3990 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1140 0.6790 1.9390 1.7870 ;
    LAYER M1 ;
      RECT 1.3830 0.6810 1.4690 0.6990 ;
      RECT 1.2310 0.6310 1.4690 0.6810 ;
      RECT 1.3830 0.6130 1.4690 0.6310 ;
      RECT 1.2310 0.6810 1.2810 0.9560 ;
      RECT 1.2310 0.5420 1.2810 0.6310 ;
      RECT 1.1910 0.9560 1.2810 1.0060 ;
      RECT 1.1910 0.4920 1.2810 0.5420 ;
      RECT 1.1910 1.0060 1.2410 1.4260 ;
      RECT 1.1910 0.1880 1.2410 0.4920 ;
      RECT 1.0790 0.6640 1.1650 0.7500 ;
      RECT 1.0790 0.7500 1.1290 1.2260 ;
      RECT 1.0790 0.6160 1.1290 0.6640 ;
      RECT 0.5830 1.2260 1.1290 1.2760 ;
      RECT 0.7350 0.5660 1.1290 0.6160 ;
      RECT 0.7350 0.2120 0.7850 0.5660 ;
      RECT 0.5830 1.2760 0.6330 1.3930 ;
      RECT 0.5830 1.1060 0.6330 1.2260 ;
      RECT 0.5830 0.0950 0.9370 0.1450 ;
      RECT 0.5830 0.1450 0.6330 0.5980 ;
      RECT 0.8870 0.1450 0.9370 0.5040 ;
      RECT 0.2790 0.5980 0.6330 0.6480 ;
      RECT 0.2790 0.1780 0.3290 0.5980 ;
    LAYER PO ;
      RECT 0.0610 0.1010 0.0910 1.4690 ;
      RECT 0.5170 0.1010 0.5470 1.5670 ;
      RECT 0.2130 0.1010 0.2430 1.4690 ;
      RECT 0.9730 0.1010 1.0030 1.4690 ;
      RECT 0.8210 0.1010 0.8510 1.4690 ;
      RECT 0.6690 0.1010 0.6990 1.4690 ;
      RECT 1.1250 0.0540 1.1550 1.6080 ;
      RECT 1.4290 0.0690 1.4590 1.6080 ;
      RECT 1.2770 0.1010 1.3070 1.4690 ;
      RECT 0.3650 0.1010 0.3950 1.4690 ;
      RECT 1.5810 0.1010 1.6110 1.4690 ;
      RECT 1.7330 0.1010 1.7630 1.4690 ;
  END
END OAI22X1_LVT

MACRO OAI22X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.976 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.9760 1.7020 ;
        RECT 0.2790 0.9580 0.3290 1.6420 ;
        RECT 1.0390 1.3630 1.0890 1.6420 ;
        RECT 0.8870 1.3350 0.9370 1.6420 ;
        RECT 1.4950 1.1330 1.5450 1.6420 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3430 0.5300 1.8360 0.5420 ;
        RECT 1.7860 0.5420 1.8360 0.9560 ;
        RECT 1.3430 0.4920 1.9110 0.5300 ;
        RECT 1.3430 0.9560 1.8360 1.0060 ;
        RECT 1.7510 0.3920 1.9110 0.4920 ;
        RECT 1.6470 0.1880 1.6970 0.4920 ;
        RECT 1.3430 0.1880 1.3930 0.4920 ;
        RECT 1.6470 1.0060 1.6970 1.4260 ;
        RECT 1.3430 1.0060 1.3930 1.4260 ;
    END
    ANTENNADIFFAREA 0.2464 ;
  END Y

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 0.8540 0.7090 0.9670 ;
        RECT 0.5600 0.9670 0.7090 0.9860 ;
        RECT 0.6590 0.7230 0.7090 0.8540 ;
    END
    ANTENNAGATEAREA 0.0276 ;
  END A4

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8110 0.7150 0.8610 1.0020 ;
        RECT 0.8110 1.0020 0.9680 1.1390 ;
    END
    ANTENNAGATEAREA 0.0276 ;
  END A3

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 1.4610 0.5730 1.5750 ;
        RECT 0.4260 1.4600 0.5730 1.4610 ;
    END
    ANTENNAGATEAREA 0.0276 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7010 0.3590 0.7100 ;
        RECT 0.2490 0.7100 0.4210 0.8150 ;
        RECT 0.2710 0.8150 0.4210 0.8170 ;
    END
    ANTENNAGATEAREA 0.0276 ;
  END A1

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.9760 0.0300 ;
        RECT 0.4310 0.0300 0.4810 0.5120 ;
        RECT 1.4950 0.0300 1.5450 0.3990 ;
        RECT 1.0390 0.0300 1.0890 0.4040 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1130 0.6790 2.0920 1.7870 ;
    LAYER M1 ;
      RECT 1.2310 0.6310 1.6210 0.6810 ;
      RECT 1.5350 0.6810 1.6210 0.6990 ;
      RECT 1.5350 0.6130 1.6210 0.6310 ;
      RECT 1.3740 0.6810 1.4600 0.6990 ;
      RECT 1.3740 0.6130 1.4600 0.6310 ;
      RECT 1.2310 0.6810 1.2810 0.9560 ;
      RECT 1.2310 0.5420 1.2810 0.6310 ;
      RECT 1.1910 0.9560 1.2810 1.0060 ;
      RECT 1.1910 0.4920 1.2810 0.5420 ;
      RECT 1.1910 1.0060 1.2410 1.4260 ;
      RECT 1.1910 0.1880 1.2410 0.4920 ;
      RECT 1.0790 0.6640 1.1650 0.7500 ;
      RECT 1.0790 0.7500 1.1290 1.2260 ;
      RECT 1.0790 0.6160 1.1290 0.6640 ;
      RECT 0.5830 1.2260 1.1290 1.2760 ;
      RECT 0.7350 0.5660 1.1290 0.6160 ;
      RECT 0.7350 0.2120 0.7850 0.5660 ;
      RECT 0.5830 1.2760 0.6330 1.3930 ;
      RECT 0.5830 1.1060 0.6330 1.2260 ;
      RECT 0.5830 0.0950 0.9370 0.1450 ;
      RECT 0.8870 0.1450 0.9370 0.5040 ;
      RECT 0.5830 0.1450 0.6330 0.5980 ;
      RECT 0.2790 0.5980 0.6330 0.6480 ;
      RECT 0.2790 0.1780 0.3290 0.5980 ;
    LAYER PO ;
      RECT 1.7330 0.1010 1.7630 1.4690 ;
      RECT 0.8210 0.1010 0.8510 1.4690 ;
      RECT 0.6690 0.1010 0.6990 1.4690 ;
      RECT 1.4290 0.0690 1.4590 1.6080 ;
      RECT 0.3650 0.1010 0.3950 1.4690 ;
      RECT 1.2770 0.1010 1.3070 1.4690 ;
      RECT 1.8850 0.1010 1.9150 1.4690 ;
      RECT 0.5170 0.1010 0.5470 1.5670 ;
      RECT 1.5810 0.0690 1.6110 1.6080 ;
      RECT 1.1250 0.0540 1.1550 1.6080 ;
      RECT 0.9730 0.1010 1.0030 1.4690 ;
      RECT 0.0610 0.1010 0.0910 1.4690 ;
      RECT 0.2130 0.1010 0.2430 1.4690 ;
  END
END OAI22X2_LVT

MACRO NOR2X0_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.52 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3130 0.4900 1.4230 0.5110 ;
        RECT 1.1910 0.4400 1.4230 0.4900 ;
        RECT 1.3450 0.5110 1.3950 0.7740 ;
        RECT 1.3130 0.4010 1.4230 0.4400 ;
        RECT 1.1910 0.4900 1.2410 0.4920 ;
        RECT 1.1910 0.1310 1.2410 0.4400 ;
        RECT 1.1910 0.7740 1.3950 0.8240 ;
        RECT 1.1910 0.8240 1.2410 1.5520 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.5200 1.7020 ;
        RECT 0.7350 0.9880 0.7850 1.6420 ;
        RECT 1.0390 0.9110 1.0890 1.6420 ;
        RECT 0.2790 0.9110 0.3290 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.5200 0.0300 ;
        RECT 0.7350 0.0300 0.7850 0.2950 ;
        RECT 1.0390 0.0300 1.0890 0.3870 ;
        RECT 0.4310 0.0300 0.4810 0.3300 ;
    END
  END VSS

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4910 0.5530 0.6650 0.7110 ;
    END
    ANTENNAGATEAREA 0.0303 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6570 0.4210 0.8510 ;
    END
    ANTENNAGATEAREA 0.0303 ;
  END A1
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.6350 1.7730 ;
    LAYER M1 ;
      RECT 0.2790 0.3830 0.7750 0.4330 ;
      RECT 0.5830 0.8130 0.7750 0.8630 ;
      RECT 0.5830 0.1740 0.6330 0.3830 ;
      RECT 0.5830 0.8630 0.6330 1.5520 ;
      RECT 0.7250 0.4330 0.7750 0.6660 ;
      RECT 0.7250 0.6660 0.8770 0.7160 ;
      RECT 0.7250 0.7160 0.7750 0.8130 ;
      RECT 0.2790 0.1740 0.3290 0.3830 ;
      RECT 1.0100 0.6610 1.1810 0.7110 ;
      RECT 0.8870 0.7730 1.0600 0.8230 ;
      RECT 1.0100 0.7110 1.0600 0.7730 ;
      RECT 1.0100 0.5520 1.0600 0.6610 ;
      RECT 0.8870 0.5020 1.0610 0.5520 ;
      RECT 0.8870 0.8230 0.9370 1.1520 ;
      RECT 0.8870 0.1310 0.9370 0.5020 ;
    LAYER PO ;
      RECT 1.1250 0.0710 1.1550 1.6120 ;
      RECT 1.2770 0.0710 1.3070 1.6120 ;
      RECT 0.8210 0.0710 0.8510 1.6120 ;
      RECT 0.9730 0.0710 1.0030 1.6120 ;
      RECT 0.0610 0.0710 0.0910 1.6120 ;
      RECT 1.4290 0.0710 1.4590 1.6120 ;
      RECT 0.2130 0.0710 0.2430 1.6120 ;
      RECT 0.6690 0.0710 0.6990 1.6120 ;
      RECT 0.3650 0.0710 0.3950 1.6120 ;
      RECT 0.5170 0.0710 0.5470 1.6120 ;
  END
END NOR2X0_LVT

MACRO NOR2X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.52 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3130 0.4900 1.4230 0.5110 ;
        RECT 1.1910 0.4400 1.4230 0.4900 ;
        RECT 1.3450 0.5110 1.3950 0.7740 ;
        RECT 1.3130 0.4010 1.4230 0.4400 ;
        RECT 1.1910 0.4900 1.2410 0.4920 ;
        RECT 1.1910 0.1310 1.2410 0.4400 ;
        RECT 1.1910 0.7740 1.3950 0.8240 ;
        RECT 1.1910 0.8240 1.2410 1.5520 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6440 1.5200 1.7000 ;
        RECT 0.7350 0.9880 0.7850 1.6440 ;
        RECT 1.0390 0.9110 1.0890 1.6440 ;
        RECT 0.2790 0.9110 0.3290 1.6440 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0280 1.5200 0.0280 ;
        RECT 0.7350 0.0280 0.7850 0.2950 ;
        RECT 1.0390 0.0280 1.0890 0.3870 ;
        RECT 0.4310 0.0280 0.4810 0.3300 ;
    END
  END VSS

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4890 0.5530 0.6630 0.7330 ;
    END
    ANTENNAGATEAREA 0.0303 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6310 0.4210 0.8150 ;
    END
    ANTENNAGATEAREA 0.0303 ;
  END A1
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.6350 1.7730 ;
    LAYER M1 ;
      RECT 0.2790 0.3830 0.7750 0.4330 ;
      RECT 0.7250 0.4330 0.7750 0.6660 ;
      RECT 0.7250 0.6660 0.8770 0.7160 ;
      RECT 0.7250 0.7160 0.7750 0.8130 ;
      RECT 0.5830 0.8130 0.7750 0.8630 ;
      RECT 0.5830 0.1740 0.6330 0.3830 ;
      RECT 0.5830 0.8630 0.6330 1.5520 ;
      RECT 0.2790 0.1740 0.3290 0.3830 ;
      RECT 1.0100 0.6610 1.1810 0.7110 ;
      RECT 0.8870 0.7730 1.0600 0.8230 ;
      RECT 1.0100 0.7110 1.0600 0.7730 ;
      RECT 1.0100 0.5520 1.0600 0.6610 ;
      RECT 0.8870 0.5020 1.0610 0.5520 ;
      RECT 0.8870 0.8230 0.9370 1.1520 ;
      RECT 0.8870 0.1310 0.9370 0.5020 ;
    LAYER PO ;
      RECT 1.1250 0.0710 1.1550 1.6120 ;
      RECT 1.2770 0.0710 1.3070 1.6120 ;
      RECT 0.8210 0.0710 0.8510 1.6120 ;
      RECT 0.9730 0.0710 1.0030 1.6120 ;
      RECT 0.0610 0.0710 0.0910 1.6120 ;
      RECT 1.4290 0.0710 1.4590 1.6120 ;
      RECT 0.2130 0.0710 0.2430 1.6120 ;
      RECT 0.6690 0.0710 0.6990 1.6120 ;
      RECT 0.3650 0.0710 0.3950 1.6120 ;
      RECT 0.5170 0.0710 0.5470 1.6120 ;
  END
END NOR2X1_LVT

MACRO NOR2X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.672 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4650 0.4010 1.5750 0.4940 ;
        RECT 1.1910 0.4940 1.5750 0.5110 ;
        RECT 1.1910 0.5110 1.5510 0.5440 ;
        RECT 1.1910 0.1310 1.2410 0.4940 ;
        RECT 1.1910 0.5440 1.2410 0.5460 ;
        RECT 1.5010 0.5440 1.5510 0.8030 ;
        RECT 1.1910 0.8030 1.5510 0.8530 ;
        RECT 1.1910 0.8530 1.2410 1.5520 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.6720 1.7020 ;
        RECT 0.7350 0.9730 0.7850 1.6420 ;
        RECT 1.3430 0.9110 1.3930 1.6420 ;
        RECT 1.0390 1.0040 1.0890 1.6420 ;
        RECT 0.2790 0.9110 0.3290 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.6720 0.0300 ;
        RECT 0.4310 0.0300 0.4810 0.3190 ;
        RECT 0.7350 0.0300 0.7850 0.3190 ;
        RECT 1.3430 0.0300 1.3930 0.3870 ;
        RECT 1.0390 0.0300 1.0890 0.3870 ;
    END
  END VSS

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4890 0.5530 0.6630 0.7330 ;
    END
    ANTENNAGATEAREA 0.03 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6310 0.4210 0.8150 ;
    END
    ANTENNAGATEAREA 0.03 ;
  END A1
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.7870 1.7730 ;
    LAYER M1 ;
      RECT 0.2790 0.3830 0.7750 0.4330 ;
      RECT 0.7250 0.4330 0.7750 0.6660 ;
      RECT 0.7250 0.6660 0.8770 0.7160 ;
      RECT 0.7250 0.7160 0.7750 0.8020 ;
      RECT 0.5830 0.8020 0.7750 0.8520 ;
      RECT 0.5830 0.1310 0.6330 0.3830 ;
      RECT 0.5830 0.8520 0.6330 1.5520 ;
      RECT 0.2790 0.1310 0.3290 0.3830 ;
      RECT 1.0100 0.6610 1.3330 0.7110 ;
      RECT 0.8870 0.1310 0.9370 0.5010 ;
      RECT 0.8870 0.8530 0.9370 1.1520 ;
      RECT 0.8870 0.7920 0.9370 0.8030 ;
      RECT 1.0100 0.5510 1.0600 0.6610 ;
      RECT 1.0100 0.7110 1.0600 0.8030 ;
      RECT 0.8870 0.5010 1.0600 0.5510 ;
      RECT 0.8870 0.8030 1.0610 0.8530 ;
    LAYER PO ;
      RECT 1.1250 0.0710 1.1550 1.6120 ;
      RECT 1.2770 0.0710 1.3070 1.6120 ;
      RECT 1.4290 0.0710 1.4590 1.6120 ;
      RECT 0.8210 0.0710 0.8510 1.6120 ;
      RECT 0.9730 0.0710 1.0030 1.6120 ;
      RECT 0.0610 0.0710 0.0910 1.6120 ;
      RECT 1.5810 0.0710 1.6110 1.6120 ;
      RECT 0.2130 0.0710 0.2430 1.6120 ;
      RECT 0.6690 0.0710 0.6990 1.6120 ;
      RECT 0.3650 0.0710 0.3950 1.6120 ;
      RECT 0.5170 0.0710 0.5470 1.6120 ;
  END
END NOR2X2_LVT

MACRO NOR2X4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.976 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7690 0.4010 1.8790 0.5010 ;
        RECT 1.1910 0.5010 1.8790 0.5110 ;
        RECT 1.1910 0.5110 1.8310 0.5510 ;
        RECT 1.4950 0.1310 1.5450 0.5010 ;
        RECT 1.1910 0.1310 1.2410 0.5010 ;
        RECT 1.4950 0.5510 1.5450 0.5530 ;
        RECT 1.1910 0.5510 1.2410 0.5530 ;
        RECT 1.7810 0.5510 1.8310 0.7760 ;
        RECT 1.1910 0.7760 1.8310 0.8260 ;
        RECT 1.4950 0.8260 1.5450 1.5340 ;
        RECT 1.1910 0.8260 1.2410 1.5340 ;
    END
    ANTENNADIFFAREA 0.2976 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.9760 1.7020 ;
        RECT 1.6470 0.9110 1.6970 1.6420 ;
        RECT 1.0390 0.9110 1.0890 1.6420 ;
        RECT 1.3430 0.9110 1.3930 1.6420 ;
        RECT 0.7350 0.9730 0.7850 1.6420 ;
        RECT 0.2790 0.9110 0.3290 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.9760 0.0300 ;
        RECT 0.7350 0.0300 0.7850 0.3190 ;
        RECT 0.4310 0.0300 0.4810 0.3460 ;
        RECT 1.6470 0.0300 1.6970 0.4110 ;
        RECT 1.0390 0.0300 1.0890 0.4110 ;
        RECT 1.3430 0.0300 1.3930 0.4110 ;
    END
  END VSS

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4890 0.5530 0.6630 0.7330 ;
    END
    ANTENNAGATEAREA 0.0288 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6310 0.4210 0.8150 ;
    END
    ANTENNAGATEAREA 0.0288 ;
  END A1
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 2.0910 1.7730 ;
    LAYER M1 ;
      RECT 0.2790 0.3970 0.7750 0.4470 ;
      RECT 0.7250 0.4470 0.7750 0.6660 ;
      RECT 0.7250 0.6660 0.8770 0.7160 ;
      RECT 0.7250 0.7160 0.7750 0.8010 ;
      RECT 0.5830 0.8010 0.7750 0.8510 ;
      RECT 0.5830 0.1750 0.6330 0.3970 ;
      RECT 0.5830 0.8510 0.6330 1.5520 ;
      RECT 0.2790 0.1750 0.3290 0.3970 ;
      RECT 1.0100 0.6610 1.6370 0.7110 ;
      RECT 0.8870 0.1310 0.9370 0.5010 ;
      RECT 0.8870 0.8250 0.9370 1.1520 ;
      RECT 1.0100 0.5510 1.0600 0.6610 ;
      RECT 1.0100 0.7110 1.0600 0.7750 ;
      RECT 0.8870 0.5010 1.0600 0.5510 ;
      RECT 0.8870 0.7750 1.0610 0.8250 ;
      RECT 1.0100 0.8250 1.0600 0.8280 ;
    LAYER PO ;
      RECT 1.4290 0.0710 1.4590 1.6120 ;
      RECT 1.2770 0.0710 1.3070 1.6120 ;
      RECT 1.1250 0.0710 1.1550 1.6120 ;
      RECT 1.5810 0.0710 1.6110 1.6120 ;
      RECT 1.7330 0.0710 1.7630 1.6120 ;
      RECT 0.8210 0.0710 0.8510 1.6120 ;
      RECT 0.9730 0.0710 1.0030 1.6120 ;
      RECT 0.0610 0.0710 0.0910 1.6120 ;
      RECT 1.8850 0.0710 1.9150 1.6120 ;
      RECT 0.2130 0.0710 0.2430 1.6120 ;
      RECT 0.6690 0.0710 0.6990 1.6120 ;
      RECT 0.3650 0.0710 0.3950 1.6120 ;
      RECT 0.5170 0.0710 0.5470 1.6120 ;
  END
END NOR2X4_LVT

MACRO NOR3X0_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.672 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4650 0.4010 1.5750 0.4370 ;
        RECT 1.3430 0.4370 1.5750 0.4870 ;
        RECT 1.4650 0.4870 1.5750 0.5110 ;
        RECT 1.3430 0.4870 1.3930 0.4890 ;
        RECT 1.3430 0.1280 1.3930 0.4370 ;
        RECT 1.4970 0.5110 1.5470 0.7630 ;
        RECT 1.3430 0.7630 1.5470 0.8130 ;
        RECT 1.3430 0.8130 1.3930 1.5490 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6630 0.4170 0.8150 ;
        RECT 0.3500 0.6450 0.4100 0.6630 ;
    END
    ANTENNAGATEAREA 0.0288 ;
  END A1

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6600 0.5530 0.8150 0.7470 ;
    END
    ANTENNAGATEAREA 0.0288 ;
  END A3

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.6720 1.7020 ;
        RECT 1.1910 1.0010 1.2410 1.6420 ;
        RECT 0.8870 0.9620 0.9370 1.6420 ;
        RECT 0.2790 0.9100 0.3290 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.6720 0.0300 ;
        RECT 0.8870 0.0300 0.9370 0.2000 ;
        RECT 0.7350 0.0300 0.7850 0.2240 ;
        RECT 0.4310 0.0300 0.4810 0.2240 ;
        RECT 1.1910 0.0300 1.2410 0.3840 ;
    END
  END VSS

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 0.4420 0.5570 0.5110 ;
        RECT 0.5070 0.5110 0.5570 0.7470 ;
        RECT 0.4010 0.4010 0.5370 0.4420 ;
    END
    ANTENNAGATEAREA 0.0288 ;
  END A2
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.7870 1.7730 ;
    LAYER M1 ;
      RECT 0.7350 0.8200 0.9310 0.8700 ;
      RECT 0.8810 0.7970 0.9310 0.8200 ;
      RECT 0.8810 0.7470 1.0290 0.7970 ;
      RECT 0.8810 0.3250 0.9310 0.7470 ;
      RECT 0.2630 0.2750 0.9310 0.3250 ;
      RECT 0.8810 0.2720 0.9310 0.2750 ;
      RECT 0.5830 0.1670 0.6330 0.2750 ;
      RECT 0.7350 0.8700 0.7850 1.5490 ;
      RECT 0.2790 0.1670 0.3290 0.2750 ;
      RECT 1.1620 0.6610 1.3330 0.7110 ;
      RECT 1.0390 0.8470 1.2120 0.8970 ;
      RECT 1.1620 0.7110 1.2120 0.8470 ;
      RECT 1.1620 0.5480 1.2120 0.6610 ;
      RECT 1.0390 0.4980 1.2130 0.5480 ;
      RECT 1.0390 0.8970 1.0890 1.2330 ;
      RECT 1.0390 0.1280 1.0890 0.4980 ;
    LAYER PO ;
      RECT 1.2770 0.0680 1.3070 1.6090 ;
      RECT 1.4290 0.0680 1.4590 1.6090 ;
      RECT 0.9730 0.0680 1.0030 1.6090 ;
      RECT 1.1250 0.0680 1.1550 1.6090 ;
      RECT 1.5810 0.0700 1.6110 1.6110 ;
      RECT 0.8210 0.0680 0.8510 1.6090 ;
      RECT 0.0610 0.0680 0.0910 1.6090 ;
      RECT 0.2130 0.0680 0.2430 1.6090 ;
      RECT 0.6690 0.0680 0.6990 1.6090 ;
      RECT 0.3650 0.0680 0.3950 1.6090 ;
      RECT 0.5170 0.0680 0.5470 1.6090 ;
  END
END NOR3X0_LVT

MACRO NOR3X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.672 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4650 0.4010 1.5750 0.4370 ;
        RECT 1.3430 0.4370 1.5750 0.4870 ;
        RECT 1.4650 0.4870 1.5750 0.5110 ;
        RECT 1.3430 0.4870 1.3930 0.4890 ;
        RECT 1.3430 0.1280 1.3930 0.4370 ;
        RECT 1.4970 0.5110 1.5470 0.7630 ;
        RECT 1.3430 0.7630 1.5470 0.8130 ;
        RECT 1.3430 0.8130 1.3930 1.5490 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6630 0.4170 0.8150 ;
        RECT 0.3500 0.6450 0.4100 0.6630 ;
    END
    ANTENNAGATEAREA 0.0288 ;
  END A1

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6600 0.5530 0.8150 0.7470 ;
    END
    ANTENNAGATEAREA 0.0288 ;
  END A3

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.6720 1.7020 ;
        RECT 1.1910 1.0010 1.2410 1.6420 ;
        RECT 0.8870 0.9620 0.9370 1.6420 ;
        RECT 0.2790 0.9100 0.3290 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.6720 0.0300 ;
        RECT 0.8870 0.0300 0.9370 0.2000 ;
        RECT 0.7350 0.0300 0.7850 0.2240 ;
        RECT 0.4310 0.0300 0.4810 0.2240 ;
        RECT 1.1910 0.0300 1.2410 0.3840 ;
    END
  END VSS

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 0.4420 0.5570 0.5110 ;
        RECT 0.5070 0.5110 0.5570 0.7470 ;
        RECT 0.4010 0.4010 0.5370 0.4420 ;
    END
    ANTENNAGATEAREA 0.0288 ;
  END A2
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.7870 1.7730 ;
    LAYER M1 ;
      RECT 0.7350 0.8200 0.9310 0.8700 ;
      RECT 0.8810 0.7970 0.9310 0.8200 ;
      RECT 0.8810 0.7470 1.0290 0.7970 ;
      RECT 0.8810 0.3250 0.9310 0.7470 ;
      RECT 0.2630 0.2750 0.9310 0.3250 ;
      RECT 0.8810 0.2720 0.9310 0.2750 ;
      RECT 0.5830 0.1670 0.6330 0.2750 ;
      RECT 0.7350 0.8700 0.7850 1.5490 ;
      RECT 0.2790 0.1670 0.3290 0.2750 ;
      RECT 1.1620 0.6610 1.3330 0.7110 ;
      RECT 1.0390 0.8470 1.2120 0.8970 ;
      RECT 1.1620 0.7110 1.2120 0.8470 ;
      RECT 1.1620 0.5480 1.2120 0.6610 ;
      RECT 1.0390 0.4980 1.2130 0.5480 ;
      RECT 1.0390 0.8970 1.0890 1.2330 ;
      RECT 1.0390 0.1280 1.0890 0.4980 ;
    LAYER PO ;
      RECT 1.2770 0.0680 1.3070 1.6090 ;
      RECT 1.4290 0.0680 1.4590 1.6090 ;
      RECT 0.9730 0.0680 1.0030 1.6090 ;
      RECT 1.1250 0.0680 1.1550 1.6090 ;
      RECT 1.5810 0.0700 1.6110 1.6110 ;
      RECT 0.8210 0.0680 0.8510 1.6090 ;
      RECT 0.0610 0.0680 0.0910 1.6090 ;
      RECT 0.2130 0.0680 0.2430 1.6090 ;
      RECT 0.6690 0.0680 0.6990 1.6090 ;
      RECT 0.3650 0.0680 0.3950 1.6090 ;
      RECT 0.5170 0.0680 0.5470 1.6090 ;
  END
END NOR3X1_LVT

MACRO NOR3X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.824 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6170 0.2490 1.7270 0.3590 ;
        RECT 1.6530 0.3590 1.7030 0.5000 ;
        RECT 1.3430 0.5000 1.7030 0.5500 ;
        RECT 1.3430 0.1310 1.3930 0.5000 ;
        RECT 1.6530 0.5500 1.7030 0.8040 ;
        RECT 1.3430 0.8040 1.7030 0.8540 ;
        RECT 1.3430 0.8030 1.3930 0.8040 ;
        RECT 1.3430 0.8540 1.3930 1.5340 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6630 0.4170 0.8150 ;
        RECT 0.3500 0.6450 0.4100 0.6630 ;
    END
    ANTENNAGATEAREA 0.0285 ;
  END A1

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6600 0.5510 0.8150 0.7270 ;
    END
    ANTENNAGATEAREA 0.0285 ;
  END A3

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.8240 1.7020 ;
        RECT 1.1910 1.0040 1.2410 1.6420 ;
        RECT 1.4950 0.9110 1.5450 1.6420 ;
        RECT 0.8870 0.9620 0.9370 1.6420 ;
        RECT 0.2790 0.9100 0.3290 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.8240 0.0300 ;
        RECT 1.4950 0.0300 1.5450 0.4110 ;
        RECT 1.1910 0.0300 1.2410 0.4110 ;
        RECT 0.8870 0.0300 0.9370 0.2000 ;
        RECT 0.7350 0.0300 0.7850 0.2240 ;
        RECT 0.4310 0.0300 0.4810 0.2240 ;
    END
  END VSS

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 0.4420 0.5570 0.5110 ;
        RECT 0.5070 0.5110 0.5570 0.7470 ;
        RECT 0.4010 0.4010 0.5370 0.4420 ;
    END
    ANTENNAGATEAREA 0.0285 ;
  END A2
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.9390 1.7730 ;
    LAYER M1 ;
      RECT 0.7350 0.8320 0.9310 0.8820 ;
      RECT 0.8810 0.7970 0.9310 0.8320 ;
      RECT 0.8810 0.7470 1.0290 0.7970 ;
      RECT 0.8810 0.3250 0.9310 0.7470 ;
      RECT 0.2630 0.2750 0.9310 0.3250 ;
      RECT 0.8810 0.2720 0.9310 0.2750 ;
      RECT 0.5830 0.1670 0.6330 0.2750 ;
      RECT 0.7350 0.8820 0.7850 1.5340 ;
      RECT 0.2790 0.1670 0.3290 0.2750 ;
      RECT 1.1620 0.6610 1.4850 0.7110 ;
      RECT 1.0390 0.8980 1.0890 1.2330 ;
      RECT 1.0390 0.1280 1.0890 0.4990 ;
      RECT 1.1620 0.7110 1.2120 0.8480 ;
      RECT 1.1620 0.5490 1.2120 0.6610 ;
      RECT 1.0390 0.8480 1.2120 0.8980 ;
      RECT 1.0390 0.4990 1.2130 0.5490 ;
    LAYER PO ;
      RECT 1.5810 0.0710 1.6110 1.6120 ;
      RECT 1.4290 0.0710 1.4590 1.6120 ;
      RECT 1.2770 0.0710 1.3070 1.6120 ;
      RECT 0.9730 0.0680 1.0030 1.6090 ;
      RECT 1.1250 0.0680 1.1550 1.6090 ;
      RECT 1.7330 0.0710 1.7630 1.6110 ;
      RECT 0.8210 0.0680 0.8510 1.6090 ;
      RECT 0.0610 0.0680 0.0910 1.6090 ;
      RECT 0.2130 0.0680 0.2430 1.6090 ;
      RECT 0.6690 0.0680 0.6990 1.6090 ;
      RECT 0.3650 0.0680 0.3950 1.6090 ;
      RECT 0.5170 0.0680 0.5470 1.6090 ;
  END
END NOR3X2_LVT

MACRO NOR3X4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.128 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9210 0.4010 2.0310 0.5070 ;
        RECT 1.3430 0.5070 2.0310 0.5110 ;
        RECT 1.3430 0.5110 1.9830 0.5570 ;
        RECT 1.6470 0.1310 1.6970 0.5070 ;
        RECT 1.3430 0.1310 1.3930 0.5070 ;
        RECT 1.6470 0.5570 1.6970 0.5590 ;
        RECT 1.3430 0.5570 1.3930 0.5590 ;
        RECT 1.9330 0.5570 1.9830 0.7770 ;
        RECT 1.3430 0.7770 1.9830 0.8270 ;
        RECT 1.6470 0.8270 1.6970 1.5340 ;
        RECT 1.3430 0.8270 1.3930 1.5340 ;
    END
    ANTENNADIFFAREA 0.2976 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6630 0.4170 0.8150 ;
        RECT 0.3500 0.6450 0.4100 0.6630 ;
    END
    ANTENNAGATEAREA 0.0282 ;
  END A1

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6600 0.5530 0.8150 0.7470 ;
    END
    ANTENNAGATEAREA 0.0282 ;
  END A3

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.1280 1.7020 ;
        RECT 1.7990 0.9110 1.8490 1.6420 ;
        RECT 1.1910 1.0040 1.2410 1.6420 ;
        RECT 0.8870 0.9620 0.9370 1.6420 ;
        RECT 1.4950 0.9110 1.5450 1.6420 ;
        RECT 0.2790 0.9100 0.3290 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.1280 0.0300 ;
        RECT 1.7990 0.0300 1.8490 0.4110 ;
        RECT 1.1910 0.0300 1.2410 0.4110 ;
        RECT 1.4950 0.0300 1.5450 0.4110 ;
        RECT 0.8870 0.0300 0.9370 0.2000 ;
        RECT 0.7350 0.0300 0.7850 0.2240 ;
        RECT 0.4310 0.0300 0.4810 0.2240 ;
    END
  END VSS

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 0.4420 0.5570 0.5110 ;
        RECT 0.5070 0.5110 0.5570 0.7470 ;
        RECT 0.4010 0.4010 0.5370 0.4420 ;
    END
    ANTENNAGATEAREA 0.0282 ;
  END A2
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 2.2430 1.7730 ;
    LAYER M1 ;
      RECT 1.1620 0.6610 1.7890 0.7110 ;
      RECT 1.0390 0.1280 1.0890 0.5010 ;
      RECT 1.0390 0.8970 1.0890 1.2330 ;
      RECT 1.1620 0.5510 1.2120 0.6610 ;
      RECT 1.1620 0.7110 1.2120 0.8470 ;
      RECT 1.0390 0.5010 1.2120 0.5510 ;
      RECT 1.0400 0.8470 1.2130 0.8720 ;
      RECT 1.0390 0.8720 1.2130 0.8970 ;
      RECT 0.7350 0.8330 0.9310 0.8830 ;
      RECT 0.8810 0.7970 0.9310 0.8330 ;
      RECT 0.8810 0.7470 1.0290 0.7970 ;
      RECT 0.8810 0.3250 0.9310 0.7470 ;
      RECT 0.2630 0.2750 0.9310 0.3250 ;
      RECT 0.8810 0.2720 0.9310 0.2750 ;
      RECT 0.5830 0.1670 0.6330 0.2750 ;
      RECT 0.7350 0.8830 0.7850 1.5340 ;
      RECT 0.2790 0.1670 0.3290 0.2750 ;
    LAYER PO ;
      RECT 1.1250 0.0710 1.1550 1.6120 ;
      RECT 1.5810 0.0710 1.6110 1.6120 ;
      RECT 1.4290 0.0710 1.4590 1.6120 ;
      RECT 1.2770 0.0710 1.3070 1.6120 ;
      RECT 1.7330 0.0710 1.7630 1.6120 ;
      RECT 1.8850 0.0710 1.9150 1.6120 ;
      RECT 0.9730 0.0680 1.0030 1.6090 ;
      RECT 2.0370 0.0710 2.0670 1.6120 ;
      RECT 0.8210 0.0680 0.8510 1.6090 ;
      RECT 0.0610 0.0680 0.0910 1.6090 ;
      RECT 0.2130 0.0680 0.2430 1.6090 ;
      RECT 0.6690 0.0680 0.6990 1.6090 ;
      RECT 0.3650 0.0680 0.3950 1.6090 ;
      RECT 0.5170 0.0680 0.5470 1.6090 ;
  END
END NOR3X4_LVT

MACRO NOR4X0_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.824 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6170 0.4010 1.7270 0.4370 ;
        RECT 1.4950 0.4370 1.7270 0.4870 ;
        RECT 1.6170 0.4870 1.7270 0.5110 ;
        RECT 1.4950 0.4870 1.5450 0.4890 ;
        RECT 1.4950 0.1280 1.5450 0.4370 ;
        RECT 1.6490 0.5110 1.6990 0.8920 ;
        RECT 1.4950 0.8920 1.6990 0.9420 ;
        RECT 1.4950 0.9420 1.5450 1.5310 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8090 0.6450 0.9670 0.8150 ;
    END
    ANTENNAGATEAREA 0.0279 ;
  END A4

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5070 0.6450 0.5570 0.8570 ;
        RECT 0.4010 0.8570 0.5570 0.9500 ;
        RECT 0.4010 0.9500 0.5110 0.9670 ;
    END
    ANTENNAGATEAREA 0.0279 ;
  END A2

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.8240 1.7020 ;
        RECT 1.3430 1.0010 1.3930 1.6420 ;
        RECT 1.0390 1.0540 1.0890 1.6420 ;
        RECT 0.2790 0.9100 0.3290 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.8240 0.0300 ;
        RECT 0.7350 0.0300 0.7850 0.3420 ;
        RECT 0.4310 0.0300 0.4810 0.3310 ;
        RECT 1.3430 0.0300 1.3930 0.3840 ;
        RECT 1.0390 0.0300 1.0890 0.2920 ;
    END
  END VSS

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.0070 0.7190 1.1190 ;
        RECT 0.6590 0.6450 0.7090 1.0070 ;
    END
    ANTENNAGATEAREA 0.0279 ;
  END A3

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.4050 0.6870 ;
        RECT 0.3550 0.6870 0.4050 0.7470 ;
    END
    ANTENNAGATEAREA 0.0279 ;
  END A1
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.9390 1.7730 ;
    LAYER M1 ;
      RECT 0.2790 0.3970 1.0830 0.4470 ;
      RECT 1.0330 0.4470 1.0830 0.7470 ;
      RECT 1.0330 0.7470 1.1810 0.7970 ;
      RECT 1.0330 0.7970 1.0830 0.9030 ;
      RECT 0.8870 0.9030 1.0830 0.9530 ;
      RECT 0.5830 0.2610 0.6330 0.3970 ;
      RECT 0.8870 0.2600 0.9370 0.3970 ;
      RECT 0.8870 0.9530 0.9370 1.5350 ;
      RECT 0.8870 0.8830 0.9370 0.9030 ;
      RECT 0.2790 0.2610 0.3290 0.3970 ;
      RECT 1.3140 0.6610 1.4850 0.7110 ;
      RECT 1.1910 0.4980 1.3650 0.5480 ;
      RECT 1.3140 0.5480 1.3640 0.6610 ;
      RECT 1.3140 0.7110 1.3640 0.8500 ;
      RECT 1.1920 0.8500 1.3650 0.8750 ;
      RECT 1.1910 0.8750 1.3650 0.9000 ;
      RECT 1.1910 0.1280 1.2410 0.4980 ;
      RECT 1.1910 0.9000 1.2410 1.2240 ;
    LAYER PO ;
      RECT 1.4290 0.0680 1.4590 1.6090 ;
      RECT 1.5810 0.0680 1.6110 1.6090 ;
      RECT 1.1250 0.0680 1.1550 1.6090 ;
      RECT 1.2770 0.0680 1.3070 1.6090 ;
      RECT 0.9730 0.0680 1.0030 1.6090 ;
      RECT 1.7330 0.0720 1.7630 1.6090 ;
      RECT 0.0610 0.0720 0.0910 1.6090 ;
      RECT 0.8210 0.0720 0.8510 1.6090 ;
      RECT 0.2130 0.0720 0.2430 1.6090 ;
      RECT 0.6690 0.0720 0.6990 1.6090 ;
      RECT 0.3650 0.0720 0.3950 1.6090 ;
      RECT 0.5170 0.0720 0.5470 1.6090 ;
  END
END NOR4X0_LVT

MACRO NOR4X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.824 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6170 0.4010 1.7270 0.4370 ;
        RECT 1.4950 0.4370 1.7270 0.4870 ;
        RECT 1.6170 0.4870 1.7270 0.5110 ;
        RECT 1.4950 0.4870 1.5450 0.4890 ;
        RECT 1.4950 0.1280 1.5450 0.4370 ;
        RECT 1.6490 0.5110 1.6990 0.8920 ;
        RECT 1.4950 0.8920 1.6990 0.9420 ;
        RECT 1.4950 0.9420 1.5450 1.5310 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8090 0.6450 0.9670 0.8150 ;
    END
    ANTENNAGATEAREA 0.0279 ;
  END A4

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5070 0.6450 0.5570 0.8570 ;
        RECT 0.4010 0.8570 0.5570 0.9500 ;
        RECT 0.4010 0.9500 0.5110 0.9670 ;
    END
    ANTENNAGATEAREA 0.0279 ;
  END A2

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.8240 1.7020 ;
        RECT 1.3430 1.0930 1.3930 1.6420 ;
        RECT 1.0390 0.9770 1.0890 1.6420 ;
        RECT 0.2790 0.9100 0.3290 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.8240 0.0300 ;
        RECT 1.3430 0.0300 1.3930 0.3960 ;
        RECT 0.7350 0.0300 0.7850 0.3420 ;
        RECT 0.4310 0.0300 0.4810 0.3310 ;
        RECT 1.0390 0.0300 1.0890 0.3030 ;
    END
  END VSS

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.0090 0.7190 1.1190 ;
        RECT 0.6590 0.6450 0.7090 1.0090 ;
    END
    ANTENNAGATEAREA 0.0279 ;
  END A3

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.4050 0.6630 ;
        RECT 0.3550 0.6630 0.4050 0.7470 ;
        RECT 0.3550 0.5510 0.4050 0.5530 ;
    END
    ANTENNAGATEAREA 0.0279 ;
  END A1
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.9390 1.7730 ;
    LAYER M1 ;
      RECT 0.2790 0.3970 1.0830 0.4470 ;
      RECT 1.0330 0.4470 1.0830 0.7470 ;
      RECT 1.0330 0.7470 1.1810 0.7970 ;
      RECT 1.0330 0.7970 1.0830 0.8720 ;
      RECT 0.8870 0.8750 1.0830 0.9220 ;
      RECT 1.0270 0.8720 1.0830 0.8750 ;
      RECT 0.5830 0.2610 0.6330 0.3970 ;
      RECT 0.8870 0.2600 0.9370 0.3970 ;
      RECT 0.8870 0.9220 0.9370 1.5350 ;
      RECT 0.2790 0.2610 0.3290 0.3970 ;
      RECT 1.3140 0.6610 1.4850 0.7110 ;
      RECT 1.1910 0.4980 1.3650 0.5480 ;
      RECT 1.3140 0.5480 1.3640 0.6610 ;
      RECT 1.3140 0.7110 1.3640 0.8510 ;
      RECT 1.1920 0.8510 1.3650 0.8760 ;
      RECT 1.1910 0.8760 1.3650 0.9010 ;
      RECT 1.1910 0.1280 1.2410 0.4980 ;
      RECT 1.1910 0.9010 1.2410 1.2240 ;
    LAYER PO ;
      RECT 1.4290 0.0680 1.4590 1.6090 ;
      RECT 1.5810 0.0680 1.6110 1.6090 ;
      RECT 1.1250 0.0680 1.1550 1.6090 ;
      RECT 1.2770 0.0680 1.3070 1.6090 ;
      RECT 0.9730 0.0680 1.0030 1.6090 ;
      RECT 1.7330 0.0720 1.7630 1.6090 ;
      RECT 0.0610 0.0720 0.0910 1.6090 ;
      RECT 0.8210 0.0720 0.8510 1.6090 ;
      RECT 0.2130 0.0720 0.2430 1.6090 ;
      RECT 0.6690 0.0720 0.6990 1.6090 ;
      RECT 0.3650 0.0720 0.3950 1.6090 ;
      RECT 0.5170 0.0720 0.5470 1.6090 ;
  END
END NOR4X1_LVT

MACRO OA21X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.52 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.5200 1.7020 ;
        RECT 0.2790 0.9580 0.3290 1.6420 ;
        RECT 0.8870 1.2430 0.9370 1.6420 ;
        RECT 1.0390 1.1330 1.0890 1.6420 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3300 0.5420 1.3800 0.9560 ;
        RECT 1.1910 0.5300 1.3800 0.5420 ;
        RECT 1.1910 0.9560 1.3800 1.0060 ;
        RECT 1.1910 0.4920 1.4390 0.5300 ;
        RECT 1.1910 1.0060 1.2410 1.4260 ;
        RECT 1.3030 0.3920 1.4390 0.4920 ;
        RECT 1.1910 0.1880 1.2410 0.4920 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 0.8530 0.8610 0.9620 ;
        RECT 0.7120 0.9620 0.8610 0.9860 ;
        RECT 0.8110 0.8070 0.8610 0.8530 ;
    END
    ANTENNAGATEAREA 0.0135 ;
  END A3

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4000 1.4610 0.5730 1.5750 ;
        RECT 0.4260 1.4600 0.5730 1.4610 ;
    END
    ANTENNAGATEAREA 0.027 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7010 0.3590 0.7170 ;
        RECT 0.2490 0.7170 0.4210 0.8100 ;
        RECT 0.2710 0.8100 0.4210 0.8170 ;
    END
    ANTENNAGATEAREA 0.027 ;
  END A1

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.5200 0.0300 ;
        RECT 0.4310 0.0300 0.4810 0.5120 ;
        RECT 1.0390 0.0300 1.0890 0.3990 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.6350 1.7870 ;
    LAYER M1 ;
      RECT 1.0790 0.6810 1.1650 0.6990 ;
      RECT 0.8870 0.6310 1.1760 0.6810 ;
      RECT 1.0790 0.6130 1.1650 0.6310 ;
      RECT 0.7350 1.1800 0.7850 1.3930 ;
      RECT 0.7350 1.1060 0.7850 1.1300 ;
      RECT 0.9130 0.6810 0.9630 1.1300 ;
      RECT 0.8870 0.1810 0.9370 0.6310 ;
      RECT 0.5830 1.1300 0.9630 1.1800 ;
      RECT 0.5830 1.1800 0.6330 1.3930 ;
      RECT 0.5830 1.1060 0.6330 1.1300 ;
      RECT 0.2790 0.5980 0.6330 0.6480 ;
      RECT 0.5830 0.4620 0.6330 0.5980 ;
      RECT 0.5830 0.4120 0.7850 0.4620 ;
      RECT 0.7350 0.1810 0.7850 0.4120 ;
      RECT 0.5830 0.1810 0.6330 0.4120 ;
      RECT 0.2790 0.1780 0.3290 0.5980 ;
    LAYER PO ;
      RECT 0.9730 0.1010 1.0030 1.4690 ;
      RECT 0.3650 0.1010 0.3950 1.4690 ;
      RECT 0.8210 0.1010 0.8510 1.4690 ;
      RECT 1.2770 0.1010 1.3070 1.4690 ;
      RECT 1.4290 0.1010 1.4590 1.4690 ;
      RECT 0.0610 0.1010 0.0910 1.4690 ;
      RECT 1.1250 0.0690 1.1550 1.6080 ;
      RECT 0.5170 0.1010 0.5470 1.5670 ;
      RECT 0.2130 0.1010 0.2430 1.4690 ;
      RECT 0.6690 0.1010 0.6990 1.4690 ;
  END
END OA21X1_LVT

MACRO OA21X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.672 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.6720 1.7020 ;
        RECT 0.2790 0.9580 0.3290 1.6420 ;
        RECT 0.8870 1.2430 0.9370 1.6420 ;
        RECT 1.1910 1.1330 1.2410 1.6420 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4820 0.5420 1.5320 0.9560 ;
        RECT 1.0390 0.5300 1.5320 0.5420 ;
        RECT 1.0390 0.9560 1.5320 1.0060 ;
        RECT 1.0390 0.4920 1.5910 0.5300 ;
        RECT 1.3430 1.0060 1.3930 1.4260 ;
        RECT 1.0390 1.0060 1.0890 1.4260 ;
        RECT 1.4550 0.3920 1.5910 0.4920 ;
        RECT 1.3430 0.1880 1.3930 0.4920 ;
        RECT 1.0390 0.1880 1.0890 0.4920 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END Y

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 0.8530 0.8610 0.9620 ;
        RECT 0.7120 0.9620 0.8610 0.9860 ;
        RECT 0.8110 0.8070 0.8610 0.8530 ;
    END
    ANTENNAGATEAREA 0.0132 ;
  END A3

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4000 1.4610 0.5730 1.5750 ;
        RECT 0.4260 1.4600 0.5730 1.4610 ;
    END
    ANTENNAGATEAREA 0.027 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7010 0.3590 0.7170 ;
        RECT 0.2490 0.7170 0.4210 0.8100 ;
        RECT 0.2710 0.8100 0.4210 0.8170 ;
    END
    ANTENNAGATEAREA 0.027 ;
  END A1

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.6720 0.0300 ;
        RECT 0.4310 0.0300 0.4810 0.5120 ;
        RECT 1.1910 0.0300 1.2410 0.3990 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.7870 1.7870 ;
    LAYER M1 ;
      RECT 1.2310 0.6810 1.3170 0.6990 ;
      RECT 0.8870 0.6310 1.3170 0.6810 ;
      RECT 1.2310 0.6130 1.3170 0.6310 ;
      RECT 1.0700 0.6810 1.1560 0.6990 ;
      RECT 1.0700 0.6130 1.1560 0.6310 ;
      RECT 0.7350 1.1800 0.7850 1.3930 ;
      RECT 0.7350 1.1060 0.7850 1.1300 ;
      RECT 0.9130 0.6810 0.9630 1.1300 ;
      RECT 0.8870 0.1810 0.9370 0.6310 ;
      RECT 0.5830 1.1300 0.9630 1.1800 ;
      RECT 0.5830 1.1800 0.6330 1.3930 ;
      RECT 0.5830 1.1060 0.6330 1.1300 ;
      RECT 0.2790 0.5980 0.6330 0.6480 ;
      RECT 0.5830 0.4620 0.6330 0.5980 ;
      RECT 0.5830 0.4120 0.7850 0.4620 ;
      RECT 0.7350 0.1810 0.7850 0.4120 ;
      RECT 0.5830 0.1810 0.6330 0.4120 ;
      RECT 0.2790 0.1780 0.3290 0.5980 ;
    LAYER PO ;
      RECT 0.9730 0.1010 1.0030 1.4690 ;
      RECT 1.1250 0.0690 1.1550 1.6080 ;
      RECT 0.3650 0.1010 0.3950 1.4690 ;
      RECT 0.8210 0.1010 0.8510 1.4690 ;
      RECT 1.4290 0.1010 1.4590 1.4690 ;
      RECT 1.5810 0.1010 1.6110 1.4690 ;
      RECT 0.0610 0.1010 0.0910 1.4690 ;
      RECT 1.2770 0.0690 1.3070 1.6080 ;
      RECT 0.5170 0.1010 0.5470 1.5670 ;
      RECT 0.2130 0.1010 0.2430 1.4690 ;
      RECT 0.6690 0.1010 0.6990 1.4690 ;
  END
END OA21X2_LVT

MACRO OA221X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.824 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7100 0.4210 0.8170 ;
        RECT 0.2490 0.7010 0.3590 0.7100 ;
    END
    ANTENNAGATEAREA 0.0228 ;
  END A1

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.8240 0.0300 ;
        RECT 1.3430 0.0300 1.3930 0.3990 ;
        RECT 0.4310 0.0300 0.4810 0.5120 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.8240 1.7020 ;
        RECT 0.2790 0.9580 0.3290 1.6420 ;
        RECT 1.3430 1.1330 1.3930 1.6420 ;
        RECT 1.0390 1.3330 1.0890 1.6420 ;
        RECT 0.8870 1.3350 0.9370 1.6420 ;
    END
  END VDD

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6590 0.7130 0.7090 0.8540 ;
        RECT 0.5530 0.8540 0.7090 0.9860 ;
    END
    ANTENNAGATEAREA 0.0228 ;
  END A4

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 1.4610 0.5730 1.5750 ;
        RECT 0.4260 1.4600 0.5730 1.4610 ;
    END
    ANTENNAGATEAREA 0.0228 ;
  END A2

  PIN A5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0230 0.5410 1.1230 0.5490 ;
        RECT 1.0090 0.5490 1.1230 0.6010 ;
        RECT 1.0090 0.6010 1.1650 0.6750 ;
        RECT 1.1150 0.6750 1.1650 0.8080 ;
    END
    ANTENNAGATEAREA 0.0174 ;
  END A5

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4950 0.5300 1.6840 0.5420 ;
        RECT 1.6340 0.5420 1.6840 0.9560 ;
        RECT 1.4950 0.4920 1.7590 0.5300 ;
        RECT 1.4950 0.9560 1.6840 1.0060 ;
        RECT 1.5990 0.3920 1.7590 0.4920 ;
        RECT 1.4950 0.1880 1.5450 0.4920 ;
        RECT 1.4950 1.0060 1.5450 1.4260 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8110 0.8420 0.8610 1.0020 ;
        RECT 0.8110 1.0020 0.9680 1.1390 ;
    END
    ANTENNAGATEAREA 0.0228 ;
  END A3
  OBS
    LAYER NWELL ;
      RECT -0.1350 0.6790 1.9400 1.7870 ;
    LAYER M1 ;
      RECT 1.3830 0.6810 1.4690 0.6990 ;
      RECT 1.2270 0.6310 1.4690 0.6810 ;
      RECT 1.3830 0.6130 1.4690 0.6310 ;
      RECT 1.2270 0.5330 1.2770 0.6310 ;
      RECT 1.2270 0.6810 1.2770 0.9030 ;
      RECT 1.1910 0.4830 1.2770 0.5330 ;
      RECT 1.0390 0.9030 1.2770 0.9530 ;
      RECT 1.1910 0.2110 1.2410 0.4830 ;
      RECT 1.1910 0.9530 1.2410 1.4270 ;
      RECT 1.0390 0.9530 1.0890 1.2130 ;
      RECT 0.5830 1.2130 1.0890 1.2630 ;
      RECT 0.5830 1.2630 0.6330 1.3930 ;
      RECT 0.5830 1.1060 0.6330 1.2130 ;
      RECT 0.2790 0.5980 0.9370 0.6480 ;
      RECT 0.8870 0.2080 0.9370 0.5980 ;
      RECT 0.5830 0.1810 0.6330 0.5980 ;
      RECT 0.2790 0.1780 0.3290 0.5980 ;
      RECT 0.7350 0.0980 1.0890 0.1480 ;
      RECT 1.0390 0.1480 1.0890 0.4310 ;
      RECT 0.7350 0.1480 0.7850 0.5010 ;
    LAYER PO ;
      RECT 1.2770 0.1010 1.3070 1.4690 ;
      RECT 0.3650 0.1010 0.3950 1.4690 ;
      RECT 0.9730 0.1010 1.0030 1.4690 ;
      RECT 0.0610 0.1010 0.0910 1.4690 ;
      RECT 1.7330 0.1010 1.7630 1.4690 ;
      RECT 1.5810 0.1010 1.6110 1.4690 ;
      RECT 1.1250 0.1010 1.1550 1.4690 ;
      RECT 1.4290 0.0690 1.4590 1.6080 ;
      RECT 0.2130 0.1010 0.2430 1.4690 ;
      RECT 0.5170 0.1010 0.5470 1.5670 ;
      RECT 0.6690 0.1010 0.6990 1.4690 ;
      RECT 0.8210 0.1010 0.8510 1.4690 ;
  END
END OA221X1_LVT

MACRO NAND3X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.672 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.6720 0.0300 ;
        RECT 0.8870 0.0300 0.9370 0.3070 ;
        RECT 1.1910 0.0300 1.2410 0.4910 ;
        RECT 0.2790 0.0300 0.3290 0.4790 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.6720 1.7020 ;
        RECT 1.1910 0.8150 1.2410 1.6420 ;
        RECT 0.2790 1.2850 0.3290 1.6420 ;
        RECT 0.5830 1.2880 0.6330 1.6420 ;
        RECT 0.8870 1.1830 0.9370 1.6420 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3430 0.8070 1.5740 0.8570 ;
        RECT 1.4640 0.8570 1.5740 0.9690 ;
        RECT 1.3430 0.8570 1.3930 1.5590 ;
        RECT 1.3830 0.5160 1.4330 0.8070 ;
        RECT 1.3430 0.4550 1.4330 0.5160 ;
        RECT 1.3430 0.1250 1.3930 0.4550 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7040 0.3590 0.7350 ;
        RECT 0.2490 0.7350 0.4210 0.7850 ;
        RECT 0.2490 0.7850 0.3590 0.8140 ;
    END
    ANTENNAGATEAREA 0.0201 ;
  END A3

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 0.7050 0.6630 0.7350 ;
        RECT 0.5530 0.7350 0.7250 0.7850 ;
        RECT 0.5530 0.7850 0.6630 0.8150 ;
    END
    ANTENNAGATEAREA 0.0201 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 1.0090 0.5110 1.0390 ;
        RECT 0.4010 1.0390 0.5730 1.0890 ;
        RECT 0.4010 1.0890 0.5110 1.1190 ;
    END
    ANTENNAGATEAREA 0.0201 ;
  END A2
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.7870 1.7730 ;
    LAYER M1 ;
      RECT 1.0790 0.6420 1.3330 0.6920 ;
      RECT 1.0790 0.5160 1.1290 0.6420 ;
      RECT 1.0790 0.6920 1.1290 0.8590 ;
      RECT 1.0390 0.4660 1.1290 0.5160 ;
      RECT 1.0390 0.8590 1.1290 0.9090 ;
      RECT 1.0390 0.1250 1.0890 0.4660 ;
      RECT 1.0390 0.9090 1.0890 1.5590 ;
      RECT 0.7770 0.7310 1.0290 0.7810 ;
      RECT 0.7770 0.6210 0.8270 0.7310 ;
      RECT 0.7770 0.7810 0.8270 1.1880 ;
      RECT 0.7350 0.5710 0.8270 0.6210 ;
      RECT 0.7350 0.1210 0.7850 0.5710 ;
      RECT 0.7350 1.2380 0.7850 1.5540 ;
      RECT 0.4310 1.1880 0.8270 1.2380 ;
      RECT 0.4310 1.2380 0.4810 1.5540 ;
    LAYER PO ;
      RECT 1.5810 0.0640 1.6110 1.6000 ;
      RECT 0.0610 0.0710 0.0910 1.6100 ;
      RECT 0.8210 0.0820 0.8510 1.6100 ;
      RECT 0.2130 0.0710 0.2430 1.6100 ;
      RECT 0.5170 0.0710 0.5470 1.6100 ;
      RECT 0.3650 0.0710 0.3950 1.6100 ;
      RECT 0.6690 0.0710 0.6990 1.6100 ;
      RECT 0.9730 0.0640 1.0030 1.6100 ;
      RECT 1.1250 0.0640 1.1550 1.6000 ;
      RECT 1.4290 0.0640 1.4590 1.6000 ;
      RECT 1.2770 0.0640 1.3070 1.6040 ;
  END
END NAND3X1_LVT

MACRO NAND3X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.824 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7350 0.4210 0.7850 ;
        RECT 0.2490 0.7040 0.3590 0.7350 ;
        RECT 0.2490 0.7850 0.3590 0.8150 ;
    END
    ANTENNAGATEAREA 0.0198 ;
  END A3

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.8240 1.7020 ;
        RECT 0.2790 1.3800 0.3290 1.6420 ;
        RECT 0.5830 1.3800 0.6330 1.6420 ;
        RECT 0.8870 1.1860 0.9370 1.6420 ;
        RECT 1.1910 0.8180 1.2410 1.6420 ;
        RECT 1.4950 0.8180 1.5450 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.8240 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.4790 ;
        RECT 1.4950 0.0300 1.5450 0.3900 ;
        RECT 1.1910 0.0300 1.2410 0.4820 ;
        RECT 0.8870 0.0300 0.9370 0.3180 ;
    END
  END VSS

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 1.0090 0.5110 1.0390 ;
        RECT 0.4010 1.0390 0.5730 1.0890 ;
        RECT 0.4010 1.0890 0.5110 1.1190 ;
    END
    ANTENNAGATEAREA 0.0198 ;
  END A2

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.5830 0.5530 1.7270 0.6630 ;
        RECT 1.5830 0.5060 1.6330 0.5530 ;
        RECT 1.5830 0.6630 1.6330 0.6920 ;
        RECT 1.3430 0.4560 1.6330 0.5060 ;
        RECT 1.3430 0.6920 1.6330 0.7420 ;
        RECT 1.3430 0.1240 1.3930 0.4560 ;
        RECT 1.3430 0.7420 1.3930 1.5590 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 0.7050 0.6630 0.7350 ;
        RECT 0.5530 0.7350 0.7250 0.7850 ;
        RECT 0.5530 0.7850 0.6630 0.8150 ;
    END
    ANTENNAGATEAREA 0.0198 ;
  END A1
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.9390 1.7730 ;
    LAYER M1 ;
      RECT 1.0790 0.5910 1.4850 0.6410 ;
      RECT 1.0790 0.6410 1.1290 0.8590 ;
      RECT 1.0790 0.5050 1.1290 0.5910 ;
      RECT 1.0390 0.8590 1.1290 0.9090 ;
      RECT 1.0390 0.4550 1.1290 0.5050 ;
      RECT 1.0390 0.9090 1.0890 1.5590 ;
      RECT 1.0390 0.1360 1.0890 0.4550 ;
      RECT 0.7770 0.7310 1.0290 0.7810 ;
      RECT 0.7770 0.6210 0.8270 0.7310 ;
      RECT 0.7770 0.7810 0.8270 1.2490 ;
      RECT 0.7350 0.5710 0.8270 0.6210 ;
      RECT 0.4310 1.2490 0.8270 1.2990 ;
      RECT 0.7350 0.1210 0.7850 0.5710 ;
      RECT 0.7350 1.2990 0.7850 1.5540 ;
      RECT 0.4310 1.2990 0.4810 1.5540 ;
    LAYER PO ;
      RECT 1.5810 0.0640 1.6110 1.6040 ;
      RECT 1.7330 0.0640 1.7630 1.6040 ;
      RECT 1.2770 0.0640 1.3070 1.6040 ;
      RECT 1.1250 0.0640 1.1550 1.6040 ;
      RECT 0.3650 0.0710 0.3950 1.6040 ;
      RECT 0.5170 0.0710 0.5470 1.6040 ;
      RECT 0.2130 0.0710 0.2430 1.6040 ;
      RECT 0.8210 0.0710 0.8510 1.6040 ;
      RECT 0.0610 0.0710 0.0910 1.6040 ;
      RECT 0.6690 0.0710 0.6990 1.6040 ;
      RECT 0.9730 0.0640 1.0030 1.6040 ;
      RECT 1.4290 0.0640 1.4590 1.6040 ;
  END
END NAND3X2_LVT

MACRO NAND3X4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.128 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7350 0.4210 0.7850 ;
        RECT 0.2490 0.7050 0.3590 0.7350 ;
        RECT 0.2490 0.7850 0.3590 0.8150 ;
    END
    ANTENNAGATEAREA 0.0198 ;
  END A3

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 0.7350 0.7250 0.7850 ;
        RECT 0.5530 0.7050 0.6630 0.7350 ;
        RECT 0.5530 0.7850 0.6630 0.8150 ;
    END
    ANTENNAGATEAREA 0.0198 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7990 0.1150 1.8490 0.5140 ;
        RECT 1.1910 0.5140 1.9540 0.5530 ;
        RECT 1.4950 0.1150 1.5450 0.5140 ;
        RECT 1.1910 0.1150 1.2410 0.5140 ;
        RECT 1.1910 0.5530 2.0410 0.5640 ;
        RECT 1.9040 0.5640 2.0410 0.6630 ;
        RECT 1.9040 0.6630 1.9540 0.7430 ;
        RECT 1.1910 0.7430 1.9540 0.7930 ;
        RECT 1.4950 0.7930 1.5450 1.5650 ;
        RECT 1.1910 0.7930 1.2410 1.5650 ;
        RECT 1.7990 0.7930 1.8490 1.5650 ;
    END
    ANTENNADIFFAREA 0.3972 ;
  END Y

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0280 2.1280 0.0280 ;
        RECT 0.8870 0.0280 0.9370 0.3310 ;
        RECT 1.6470 0.0280 1.6970 0.4130 ;
        RECT 1.3430 0.0280 1.3930 0.4130 ;
        RECT 0.2790 0.0280 0.3290 0.4790 ;
    END
  END VSS

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 1.0090 0.5110 1.0390 ;
        RECT 0.4010 1.0390 0.5730 1.0890 ;
        RECT 0.4010 1.0890 0.5110 1.1190 ;
    END
    ANTENNAGATEAREA 0.0198 ;
  END A2

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6440 2.1280 1.7000 ;
        RECT 1.3430 0.8470 1.3930 1.6440 ;
        RECT 1.6470 0.8470 1.6970 1.6440 ;
        RECT 0.8870 1.1830 0.9370 1.6440 ;
        RECT 0.2790 1.3770 0.3290 1.6440 ;
        RECT 0.5830 1.3770 0.6330 1.6440 ;
    END
  END VDD
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 2.2430 1.7730 ;
    LAYER M1 ;
      RECT 1.0790 0.6420 1.7890 0.6920 ;
      RECT 1.0790 0.5050 1.1290 0.6420 ;
      RECT 1.0790 0.6920 1.1290 0.8560 ;
      RECT 1.0390 0.4550 1.1290 0.5050 ;
      RECT 1.0390 0.8560 1.1290 0.9060 ;
      RECT 1.0390 0.1490 1.0890 0.4550 ;
      RECT 1.0390 0.9060 1.0890 1.5560 ;
      RECT 0.7770 0.7310 1.0290 0.7810 ;
      RECT 0.4310 1.2350 0.4810 1.5510 ;
      RECT 0.7770 0.6210 0.8270 0.7310 ;
      RECT 0.7770 0.7810 0.8270 1.1850 ;
      RECT 0.7350 0.5710 0.8270 0.6210 ;
      RECT 0.4310 1.1850 0.8270 1.2350 ;
      RECT 0.7350 0.1210 0.7850 0.5710 ;
      RECT 0.7350 1.2350 0.7850 1.5510 ;
    LAYER PO ;
      RECT 0.6690 0.0710 0.6990 1.6100 ;
      RECT 0.9730 0.0640 1.0030 1.6100 ;
      RECT 0.2130 0.0710 0.2430 1.6100 ;
      RECT 0.5170 0.0710 0.5470 1.6100 ;
      RECT 0.3650 0.0710 0.3950 1.6100 ;
      RECT 1.1250 0.0640 1.1550 1.6000 ;
      RECT 0.0610 0.0710 0.0910 1.6100 ;
      RECT 0.8210 0.0710 0.8510 1.6100 ;
      RECT 1.4290 0.0720 1.4590 1.6100 ;
      RECT 1.5810 0.0720 1.6110 1.6100 ;
      RECT 1.7330 0.0720 1.7630 1.6100 ;
      RECT 2.0370 0.0720 2.0670 1.6100 ;
      RECT 1.8850 0.0720 1.9150 1.6100 ;
      RECT 1.2770 0.0720 1.3070 1.6100 ;
  END
END NAND3X4_LVT

MACRO NAND4X0_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.216 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 0.7350 0.7250 0.7850 ;
        RECT 0.5530 0.7050 0.6630 0.7350 ;
        RECT 0.5530 0.7850 0.6630 0.8150 ;
    END
    ANTENNAGATEAREA 0.0276 ;
  END A2

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7350 0.4210 0.7850 ;
        RECT 0.2490 0.7050 0.3590 0.7350 ;
        RECT 0.2490 0.7850 0.3590 0.8150 ;
    END
    ANTENNAGATEAREA 0.0276 ;
  END A4

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.2160 1.7020 ;
        RECT 0.7350 1.1930 0.7850 1.6420 ;
        RECT 0.4310 1.1930 0.4810 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.2160 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.5710 ;
    END
  END VSS

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 0.8570 0.5110 0.8870 ;
        RECT 0.4010 0.8870 0.5730 0.9370 ;
        RECT 0.4010 0.9370 0.5110 0.9670 ;
    END
    ANTENNAGATEAREA 0.0276 ;
  END A3

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2790 1.0530 0.9770 1.1030 ;
        RECT 0.8870 1.1030 0.9370 1.5510 ;
        RECT 0.5830 1.1030 0.6330 1.5510 ;
        RECT 0.2790 1.1030 0.3290 1.5510 ;
        RECT 0.9270 0.8150 0.9770 1.0530 ;
        RECT 0.8570 0.7050 0.9770 0.8150 ;
        RECT 0.9270 0.6510 0.9770 0.7050 ;
        RECT 0.8870 0.6010 0.9770 0.6510 ;
        RECT 0.8870 0.1210 0.9370 0.6010 ;
    END
    ANTENNADIFFAREA 0.1834 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 0.8570 0.8150 0.8870 ;
        RECT 0.7050 0.8870 0.8770 0.9370 ;
        RECT 0.7050 0.9370 0.8150 0.9670 ;
    END
    ANTENNAGATEAREA 0.0276 ;
  END A1
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.7160 1.3310 1.7730 ;
      RECT -0.1150 0.6790 0.1910 0.7160 ;
      RECT 1.0180 0.6790 1.3310 0.7160 ;
    LAYER PO ;
      RECT 1.1250 0.0710 1.1550 1.6100 ;
      RECT 0.9730 0.0710 1.0030 1.6100 ;
      RECT 0.6690 0.0710 0.6990 1.6100 ;
      RECT 0.3650 0.0710 0.3950 1.6100 ;
      RECT 0.5170 0.0710 0.5470 1.6100 ;
      RECT 0.2130 0.0710 0.2430 1.6100 ;
      RECT 0.8210 0.0710 0.8510 1.6100 ;
      RECT 0.0610 0.0710 0.0910 1.6100 ;
  END
END NAND4X0_LVT

MACRO NAND4X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.824 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.5900 0.7050 1.7270 0.8150 ;
        RECT 1.5900 0.5640 1.6400 0.7050 ;
        RECT 1.5900 0.8150 1.6400 0.8260 ;
        RECT 1.3430 0.5140 1.6400 0.5640 ;
        RECT 1.3430 0.8260 1.6400 0.8760 ;
        RECT 1.3430 0.1150 1.3930 0.5140 ;
        RECT 1.3430 0.8760 1.3930 1.5610 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.8240 0.0300 ;
        RECT 1.0390 0.0300 1.0890 0.3220 ;
        RECT 0.2790 0.0300 0.3290 0.4790 ;
        RECT 1.4950 0.0300 1.5450 0.4130 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.8240 1.7020 ;
        RECT 1.4950 1.0040 1.5450 1.6420 ;
        RECT 0.7350 1.3770 0.7850 1.6420 ;
        RECT 0.4310 1.3770 0.4810 1.6420 ;
        RECT 1.0390 1.1830 1.0890 1.6420 ;
    END
  END VDD

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 0.7050 0.6630 0.7350 ;
        RECT 0.5530 0.7350 0.7250 0.7850 ;
        RECT 0.5530 0.7850 0.6630 0.8150 ;
    END
    ANTENNAGATEAREA 0.0183 ;
  END A2

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7050 0.3590 0.7350 ;
        RECT 0.2490 0.7350 0.4210 0.7850 ;
        RECT 0.2490 0.7850 0.3590 0.8150 ;
    END
    ANTENNAGATEAREA 0.0183 ;
  END A4

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 1.0090 0.5110 1.0390 ;
        RECT 0.4010 1.0390 0.5730 1.0890 ;
        RECT 0.4010 1.0890 0.5110 1.1190 ;
    END
    ANTENNAGATEAREA 0.0183 ;
  END A3

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 1.0090 0.8150 1.0390 ;
        RECT 0.7050 1.0390 0.8770 1.0890 ;
        RECT 0.7050 1.0890 0.8150 1.1190 ;
    END
    ANTENNAGATEAREA 0.0183 ;
  END A1
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.9390 1.7730 ;
    LAYER M1 ;
      RECT 0.9270 0.7370 1.1810 0.7870 ;
      RECT 0.9270 0.6370 0.9770 0.7370 ;
      RECT 0.8870 0.5870 0.9770 0.6370 ;
      RECT 0.8870 1.3270 0.9370 1.5510 ;
      RECT 0.8870 0.1210 0.9370 0.5870 ;
      RECT 0.2790 1.2770 0.9770 1.3270 ;
      RECT 0.9270 0.7870 0.9770 1.2770 ;
      RECT 0.5830 1.3270 0.6330 1.5510 ;
      RECT 0.2790 1.3270 0.3290 1.5510 ;
      RECT 1.2310 0.6140 1.4850 0.6640 ;
      RECT 1.2310 0.6640 1.2810 0.8560 ;
      RECT 1.2310 0.5050 1.2810 0.6140 ;
      RECT 1.1910 0.8560 1.2810 0.9060 ;
      RECT 1.1910 0.4550 1.2810 0.5050 ;
      RECT 1.1910 0.9060 1.2410 1.5560 ;
      RECT 1.1910 0.1400 1.2410 0.4550 ;
    LAYER PO ;
      RECT 0.3650 0.0710 0.3950 1.6100 ;
      RECT 0.5170 0.0710 0.5470 1.6100 ;
      RECT 0.6690 0.0710 0.6990 1.6100 ;
      RECT 0.2130 0.0710 0.2430 1.6100 ;
      RECT 1.2770 0.0640 1.3070 1.6000 ;
      RECT 1.1250 0.0640 1.1550 1.6100 ;
      RECT 0.8210 0.0710 0.8510 1.6100 ;
      RECT 1.5810 0.0710 1.6110 1.6100 ;
      RECT 0.0610 0.0710 0.0910 1.6100 ;
      RECT 1.4290 0.0720 1.4590 1.6100 ;
      RECT 0.9730 0.0710 1.0030 1.6100 ;
      RECT 1.7330 0.0640 1.7630 1.6000 ;
  END
END NAND4X1_LVT

MACRO NBUFFX16_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.648 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6600 0.7400 0.7100 ;
        RECT 0.2490 0.7100 0.3620 0.8150 ;
    END
    ANTENNAGATEAREA 0.1098 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.6480 1.7020 ;
        RECT 0.4310 0.9920 0.4810 1.6420 ;
        RECT 3.1670 0.9920 3.2170 1.6420 ;
        RECT 0.7350 0.9920 0.7850 1.6420 ;
        RECT 2.8630 0.9920 2.9130 1.6420 ;
        RECT 2.5590 0.9920 2.6090 1.6420 ;
        RECT 2.2550 0.9920 2.3050 1.6420 ;
        RECT 1.6470 0.9920 1.6970 1.6420 ;
        RECT 1.9510 0.9920 2.0010 1.6420 ;
        RECT 1.3430 0.9920 1.3930 1.6420 ;
        RECT 1.0390 0.9920 1.0890 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.6480 0.0300 ;
        RECT 0.4310 0.0300 0.4810 0.4100 ;
        RECT 3.1670 0.0300 3.2170 0.4100 ;
        RECT 2.8630 0.0300 2.9130 0.4100 ;
        RECT 0.7350 0.0300 0.7850 0.4100 ;
        RECT 2.5590 0.0300 2.6090 0.4100 ;
        RECT 2.2550 0.0300 2.3050 0.4100 ;
        RECT 1.6470 0.0300 1.6970 0.4100 ;
        RECT 1.9510 0.0300 2.0010 0.4100 ;
        RECT 1.3430 0.0300 1.3930 0.4100 ;
        RECT 1.0390 0.0300 1.0890 0.4100 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8870 0.5370 3.5510 0.5870 ;
        RECT 3.3780 0.5870 3.5510 0.6630 ;
        RECT 3.3190 0.1160 3.3690 0.5370 ;
        RECT 3.0150 0.1160 3.0650 0.5370 ;
        RECT 1.7990 0.1160 1.8490 0.5370 ;
        RECT 2.1030 0.1170 2.1530 0.5370 ;
        RECT 2.4070 0.1160 2.4570 0.5370 ;
        RECT 2.7110 0.1160 2.7610 0.5370 ;
        RECT 1.4950 0.1160 1.5450 0.5370 ;
        RECT 0.8870 0.1160 0.9370 0.5370 ;
        RECT 1.1910 0.1160 1.2410 0.5370 ;
        RECT 3.3780 0.6630 3.4280 0.8920 ;
        RECT 0.8870 0.8920 3.4280 0.9420 ;
        RECT 3.3190 0.9420 3.3690 1.5640 ;
        RECT 3.0150 0.9420 3.0650 1.5640 ;
        RECT 2.7110 0.9420 2.7610 1.5640 ;
        RECT 1.7990 0.9420 1.8490 1.5640 ;
        RECT 2.1030 0.9420 2.1530 1.5650 ;
        RECT 2.4070 0.9420 2.4570 1.5640 ;
        RECT 0.8870 0.9420 0.9370 1.5640 ;
        RECT 1.1910 0.9420 1.2410 1.5640 ;
        RECT 1.4950 0.9420 1.5450 1.5640 ;
    END
    ANTENNADIFFAREA 1.2904 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 3.7630 1.7730 ;
    LAYER M1 ;
      RECT 0.7900 0.6600 3.3240 0.7100 ;
      RECT 0.2790 0.8920 0.3290 1.5640 ;
      RECT 0.2790 0.5020 0.3290 0.5370 ;
      RECT 0.2790 0.1160 0.3290 0.5760 ;
      RECT 0.5830 0.8920 0.6330 1.5640 ;
      RECT 0.5830 0.1160 0.6330 0.5560 ;
      RECT 0.2790 0.8920 0.8360 0.9310 ;
      RECT 0.7860 0.8420 0.8360 0.9420 ;
      RECT 0.3290 0.9310 0.8360 0.9420 ;
      RECT 0.7900 0.7100 0.8400 0.8420 ;
      RECT 0.7900 0.8420 0.8370 0.8740 ;
      RECT 0.7900 0.6370 0.8400 0.6600 ;
      RECT 0.7900 0.6100 0.8370 0.6370 ;
      RECT 0.2790 0.5370 0.8370 0.5870 ;
      RECT 0.7870 0.5870 0.8370 0.6100 ;
    LAYER PO ;
      RECT 0.8210 0.0690 0.8510 1.6060 ;
      RECT 0.9730 0.0690 1.0030 1.6060 ;
      RECT 1.4290 0.0690 1.4590 1.6060 ;
      RECT 1.2770 0.0690 1.3070 1.6060 ;
      RECT 1.1250 0.0690 1.1550 1.6060 ;
      RECT 0.0610 0.0710 0.0910 1.6060 ;
      RECT 0.5170 0.0690 0.5470 1.6060 ;
      RECT 0.6690 0.0690 0.6990 1.6060 ;
      RECT 0.3650 0.0690 0.3950 1.6060 ;
      RECT 0.2130 0.0710 0.2430 1.6060 ;
      RECT 3.4050 0.0690 3.4350 1.6060 ;
      RECT 3.5570 0.0690 3.5870 1.6060 ;
      RECT 3.2530 0.0690 3.2830 1.6060 ;
      RECT 2.0370 0.0690 2.0670 1.6060 ;
      RECT 2.1890 0.0690 2.2190 1.6060 ;
      RECT 2.3410 0.0690 2.3710 1.6060 ;
      RECT 2.9490 0.0690 2.9790 1.6060 ;
      RECT 2.7970 0.0690 2.8270 1.6060 ;
      RECT 2.6450 0.0690 2.6750 1.6060 ;
      RECT 2.4930 0.0690 2.5230 1.6060 ;
      RECT 3.1010 0.0690 3.1310 1.6060 ;
      RECT 1.8850 0.0690 1.9150 1.6060 ;
      RECT 1.7330 0.0690 1.7630 1.6060 ;
      RECT 1.5810 0.0690 1.6110 1.6060 ;
  END
END NBUFFX16_LVT

MACRO NBUFFX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.216 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6750 0.4210 0.7250 ;
        RECT 0.2490 0.7250 0.3620 0.8150 ;
    END
    ANTENNAGATEAREA 0.0237 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.2160 1.7020 ;
        RECT 0.2790 0.9100 0.3290 1.6420 ;
        RECT 0.7350 0.9920 0.7850 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.2160 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.5670 ;
        RECT 0.7350 0.0300 0.7850 0.4100 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5830 0.1160 0.6330 0.5370 ;
        RECT 0.5830 0.5370 1.1190 0.5870 ;
        RECT 0.9430 0.5870 1.1190 0.6630 ;
        RECT 0.8870 0.1160 0.9370 0.5370 ;
        RECT 0.9430 0.6630 0.9930 0.8920 ;
        RECT 0.5830 0.8920 0.9930 0.9420 ;
        RECT 0.8870 0.9420 0.9370 1.5640 ;
        RECT 0.5830 0.9420 0.6330 1.5640 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.3310 1.7730 ;
    LAYER M1 ;
      RECT 0.4710 0.6600 0.8920 0.7100 ;
      RECT 0.4560 0.8870 0.5210 0.9370 ;
      RECT 0.4310 0.8870 0.4810 1.2680 ;
      RECT 0.4310 0.8870 0.4740 0.9370 ;
      RECT 0.4310 0.3000 0.4810 0.5710 ;
      RECT 0.4310 0.5320 0.5090 0.5820 ;
      RECT 0.4310 0.4970 0.4810 0.5320 ;
      RECT 0.4710 0.5320 0.5210 0.9370 ;
    LAYER PO ;
      RECT 0.0610 0.0710 0.0910 1.6060 ;
      RECT 0.3650 0.0690 0.3950 1.6060 ;
      RECT 0.2130 0.0710 0.2430 1.6060 ;
      RECT 0.5170 0.0710 0.5470 1.6060 ;
      RECT 0.6690 0.0690 0.6990 1.6060 ;
      RECT 1.1250 0.0710 1.1550 1.6060 ;
      RECT 0.9730 0.0710 1.0030 1.6060 ;
      RECT 0.8210 0.0690 0.8510 1.6060 ;
  END
END NBUFFX2_LVT

MACRO NBUFFX32_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.384 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6600 1.0440 0.7100 ;
        RECT 0.2490 0.7100 0.3620 0.8150 ;
    END
    ANTENNAGATEAREA 0.183 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 6.3840 1.7020 ;
        RECT 1.6470 0.9920 1.6970 1.6420 ;
        RECT 1.3430 0.9920 1.3930 1.6420 ;
        RECT 0.4310 0.9920 0.4810 1.6420 ;
        RECT 0.7350 0.9920 0.7850 1.6420 ;
        RECT 1.0390 0.9920 1.0890 1.6420 ;
        RECT 5.9030 0.9920 5.9530 1.6420 ;
        RECT 5.5990 0.9920 5.6490 1.6420 ;
        RECT 5.2950 0.9920 5.3450 1.6420 ;
        RECT 4.9910 0.9920 5.0410 1.6420 ;
        RECT 4.6870 0.9920 4.7370 1.6420 ;
        RECT 4.3830 0.9920 4.4330 1.6420 ;
        RECT 4.0790 0.9920 4.1290 1.6420 ;
        RECT 3.7750 0.9920 3.8250 1.6420 ;
        RECT 3.4710 0.9920 3.5210 1.6420 ;
        RECT 3.1670 0.9920 3.2170 1.6420 ;
        RECT 2.8630 0.9920 2.9130 1.6420 ;
        RECT 2.5590 0.9920 2.6090 1.6420 ;
        RECT 1.9510 0.9920 2.0010 1.6420 ;
        RECT 2.2550 0.9920 2.3050 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 6.3840 0.0300 ;
        RECT 1.6470 0.0300 1.6970 0.4100 ;
        RECT 1.3430 0.0300 1.3930 0.4100 ;
        RECT 0.4310 0.0300 0.4810 0.4100 ;
        RECT 0.7350 0.0300 0.7850 0.4100 ;
        RECT 1.0390 0.0300 1.0890 0.4100 ;
        RECT 5.9030 0.0300 5.9530 0.4100 ;
        RECT 5.5990 0.0300 5.6490 0.4100 ;
        RECT 5.2950 0.0300 5.3450 0.4100 ;
        RECT 4.9910 0.0300 5.0410 0.4100 ;
        RECT 4.6870 0.0300 4.7370 0.4100 ;
        RECT 4.3830 0.0300 4.4330 0.4100 ;
        RECT 4.0790 0.0300 4.1290 0.4100 ;
        RECT 3.7750 0.0300 3.8250 0.4100 ;
        RECT 3.4710 0.0300 3.5210 0.4100 ;
        RECT 3.1670 0.0300 3.2170 0.4100 ;
        RECT 2.8630 0.0300 2.9130 0.4100 ;
        RECT 2.5590 0.0300 2.6090 0.4100 ;
        RECT 1.9510 0.0300 2.0010 0.4100 ;
        RECT 2.2550 0.0300 2.3050 0.4100 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.9270 0.9420 3.9770 1.5640 ;
        RECT 4.2310 0.9420 4.2810 1.5640 ;
        RECT 4.5350 0.9420 4.5850 1.5640 ;
        RECT 4.8390 0.9420 4.8890 1.5640 ;
        RECT 5.1430 0.9420 5.1930 1.5640 ;
        RECT 5.4470 0.9420 5.4970 1.5640 ;
        RECT 5.7510 0.9420 5.8010 1.5640 ;
        RECT 6.0550 0.9420 6.1050 1.5640 ;
        RECT 2.4070 0.9420 2.4570 1.5650 ;
        RECT 2.7110 0.9420 2.7610 1.5640 ;
        RECT 2.1030 0.9420 2.1530 1.5640 ;
        RECT 3.0150 0.9420 3.0650 1.5640 ;
        RECT 3.3190 0.9420 3.3690 1.5640 ;
        RECT 3.6230 0.9420 3.6730 1.5640 ;
        RECT 1.7990 0.9420 1.8490 1.5640 ;
        RECT 1.4950 0.9420 1.5450 1.5640 ;
        RECT 1.1910 0.9420 1.2410 1.5640 ;
        RECT 1.1910 0.8920 6.1640 0.9420 ;
        RECT 6.1140 0.6630 6.1640 0.8920 ;
        RECT 1.1910 0.5370 6.2870 0.5870 ;
        RECT 1.7990 0.1160 1.8490 0.5370 ;
        RECT 3.0150 0.1160 3.0650 0.5370 ;
        RECT 2.7110 0.1160 2.7610 0.5370 ;
        RECT 2.4070 0.1170 2.4570 0.5370 ;
        RECT 2.1030 0.1160 2.1530 0.5370 ;
        RECT 3.3190 0.1160 3.3690 0.5370 ;
        RECT 3.6230 0.1160 3.6730 0.5370 ;
        RECT 1.4950 0.1160 1.5450 0.5370 ;
        RECT 1.1910 0.1160 1.2410 0.5370 ;
        RECT 6.1140 0.5870 6.2870 0.6630 ;
        RECT 3.9270 0.1160 3.9770 0.5370 ;
        RECT 4.2310 0.1160 4.2810 0.5370 ;
        RECT 4.5350 0.1160 4.5850 0.5370 ;
        RECT 4.8390 0.1160 4.8890 0.5370 ;
        RECT 5.1430 0.1160 5.1930 0.5370 ;
        RECT 5.4470 0.1160 5.4970 0.5370 ;
        RECT 5.7510 0.1160 5.8010 0.5370 ;
        RECT 6.0550 0.1160 6.1050 0.5370 ;
    END
    ANTENNADIFFAREA 2.4808 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 6.4990 1.7730 ;
    LAYER M1 ;
      RECT 1.0940 0.6600 6.0600 0.7100 ;
      RECT 0.2790 0.8920 0.3290 1.5640 ;
      RECT 0.2790 0.5020 0.3290 0.5370 ;
      RECT 0.2790 0.1160 0.3290 0.5760 ;
      RECT 0.5830 0.8920 0.6330 1.5640 ;
      RECT 0.5830 0.1160 0.6330 0.5760 ;
      RECT 0.8870 0.8920 0.9370 1.5640 ;
      RECT 0.8870 0.1160 0.9370 0.5760 ;
      RECT 0.2790 0.8920 1.1410 0.9310 ;
      RECT 0.3290 0.9310 1.1410 0.9420 ;
      RECT 1.0940 0.7100 1.1440 0.8180 ;
      RECT 1.0910 0.8180 1.1440 0.8420 ;
      RECT 1.0910 0.8420 1.1410 0.8920 ;
      RECT 1.0940 0.6370 1.1440 0.6600 ;
      RECT 1.0940 0.6100 1.1410 0.6370 ;
      RECT 0.2790 0.5370 1.1410 0.5870 ;
      RECT 1.0910 0.5870 1.1410 0.6100 ;
    LAYER PO ;
      RECT 2.7970 0.0690 2.8270 1.6060 ;
      RECT 3.4050 0.0690 3.4350 1.6060 ;
      RECT 2.1890 0.0690 2.2190 1.6060 ;
      RECT 2.0370 0.0690 2.0670 1.6060 ;
      RECT 1.8850 0.0690 1.9150 1.6060 ;
      RECT 1.1250 0.0690 1.1550 1.6060 ;
      RECT 1.2770 0.0690 1.3070 1.6060 ;
      RECT 1.7330 0.0690 1.7630 1.6060 ;
      RECT 1.5810 0.0690 1.6110 1.6060 ;
      RECT 1.4290 0.0690 1.4590 1.6060 ;
      RECT 0.0610 0.0690 0.0910 1.6060 ;
      RECT 0.5170 0.0690 0.5470 1.6060 ;
      RECT 0.6690 0.0690 0.6990 1.6060 ;
      RECT 0.8210 0.0690 0.8510 1.6060 ;
      RECT 0.3650 0.0690 0.3950 1.6060 ;
      RECT 0.2130 0.0690 0.2430 1.6060 ;
      RECT 0.9730 0.0690 1.0030 1.6060 ;
      RECT 6.2930 0.0690 6.3230 1.6060 ;
      RECT 6.1410 0.0690 6.1710 1.6060 ;
      RECT 5.9890 0.0690 6.0190 1.6060 ;
      RECT 5.8370 0.0690 5.8670 1.6060 ;
      RECT 5.5330 0.0690 5.5630 1.6060 ;
      RECT 5.6850 0.0690 5.7150 1.6060 ;
      RECT 5.2290 0.0690 5.2590 1.6060 ;
      RECT 5.3810 0.0690 5.4110 1.6060 ;
      RECT 5.0770 0.0690 5.1070 1.6060 ;
      RECT 4.9250 0.0690 4.9550 1.6060 ;
      RECT 4.7730 0.0690 4.8030 1.6060 ;
      RECT 4.6210 0.0690 4.6510 1.6060 ;
      RECT 4.3170 0.0690 4.3470 1.6060 ;
      RECT 4.4690 0.0690 4.4990 1.6060 ;
      RECT 3.7090 0.0690 3.7390 1.6060 ;
      RECT 3.8610 0.0690 3.8910 1.6060 ;
      RECT 3.5570 0.0690 3.5870 1.6060 ;
      RECT 4.0130 0.0690 4.0430 1.6060 ;
      RECT 4.1650 0.0690 4.1950 1.6060 ;
      RECT 2.3410 0.0690 2.3710 1.6060 ;
      RECT 2.4930 0.0690 2.5230 1.6060 ;
      RECT 2.6450 0.0690 2.6750 1.6060 ;
      RECT 3.2530 0.0690 3.2830 1.6060 ;
      RECT 3.1010 0.0690 3.1310 1.6060 ;
      RECT 2.9490 0.0690 2.9790 1.6060 ;
  END
END NBUFFX32_LVT

MACRO NBUFFX4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.52 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6550 0.4360 0.7050 ;
        RECT 0.2490 0.7050 0.3620 0.8150 ;
    END
    ANTENNAGATEAREA 0.0366 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.5200 1.7020 ;
        RECT 0.2790 0.9870 0.3290 1.6420 ;
        RECT 1.0390 0.9920 1.0890 1.6420 ;
        RECT 0.7350 0.9920 0.7850 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.5200 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.4050 ;
        RECT 1.0390 0.0300 1.0890 0.4100 ;
        RECT 0.7350 0.0300 0.7850 0.4100 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5830 0.5370 1.4230 0.5870 ;
        RECT 1.2460 0.5870 1.4230 0.6630 ;
        RECT 1.1910 0.1160 1.2410 0.5370 ;
        RECT 0.5830 0.1160 0.6330 0.5370 ;
        RECT 0.8870 0.1160 0.9370 0.5370 ;
        RECT 1.2460 0.6630 1.2960 0.8920 ;
        RECT 0.5830 0.8920 1.2960 0.9420 ;
        RECT 0.5830 0.9420 0.6330 1.5640 ;
        RECT 0.8870 0.9420 0.9370 1.5640 ;
        RECT 1.1910 0.9420 1.2410 1.5640 ;
    END
    ANTENNADIFFAREA 0.3976 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1120 0.6790 1.6350 1.7730 ;
    LAYER M1 ;
      RECT 0.4870 0.6600 1.1960 0.7100 ;
      RECT 0.4310 0.8220 0.4810 1.5590 ;
      RECT 0.4310 0.5320 0.5210 0.5820 ;
      RECT 0.4310 0.8870 0.4740 0.9370 ;
      RECT 0.4310 0.4970 0.4810 0.5320 ;
      RECT 0.4310 0.1110 0.4810 0.5710 ;
      RECT 0.4560 0.8220 0.5370 0.8420 ;
      RECT 0.4560 0.8420 0.5330 0.8720 ;
      RECT 0.4870 0.6370 0.5370 0.8220 ;
      RECT 0.4830 0.5320 0.5330 0.6050 ;
      RECT 0.4860 0.6050 0.5330 0.6370 ;
    LAYER PO ;
      RECT 0.0610 0.0710 0.0910 1.6060 ;
      RECT 0.3650 0.0690 0.3950 1.6060 ;
      RECT 0.2130 0.0710 0.2430 1.6060 ;
      RECT 1.4290 0.0650 1.4590 1.6000 ;
      RECT 1.2770 0.0650 1.3070 1.6000 ;
      RECT 0.5170 0.0710 0.5470 1.6060 ;
      RECT 0.6690 0.0690 0.6990 1.6060 ;
      RECT 1.1250 0.0690 1.1550 1.6060 ;
      RECT 0.9730 0.0690 1.0030 1.6060 ;
      RECT 0.8210 0.0690 0.8510 1.6060 ;
  END
END NBUFFX4_LVT

MACRO NBUFFX8_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.28 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6600 0.5880 0.7100 ;
        RECT 0.2490 0.7100 0.3620 0.8150 ;
    END
    ANTENNAGATEAREA 0.0732 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.2800 1.7020 ;
        RECT 0.4310 0.9920 0.4810 1.6420 ;
        RECT 1.4950 0.9920 1.5450 1.6420 ;
        RECT 1.7990 0.9920 1.8490 1.6420 ;
        RECT 1.1910 0.9920 1.2410 1.6420 ;
        RECT 0.8870 0.9920 0.9370 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.2800 0.0300 ;
        RECT 0.4310 0.0300 0.4810 0.4100 ;
        RECT 1.4950 0.0300 1.5450 0.4100 ;
        RECT 1.7990 0.0300 1.8490 0.4100 ;
        RECT 1.1910 0.0300 1.2410 0.4100 ;
        RECT 0.8870 0.0300 0.9370 0.4100 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7350 0.5370 2.1830 0.5870 ;
        RECT 2.0070 0.5870 2.1830 0.6630 ;
        RECT 1.6470 0.1160 1.6970 0.5370 ;
        RECT 1.9510 0.1170 2.0010 0.5370 ;
        RECT 1.3430 0.1160 1.3930 0.5370 ;
        RECT 0.7350 0.1160 0.7850 0.5370 ;
        RECT 1.0390 0.1160 1.0890 0.5370 ;
        RECT 2.0070 0.6630 2.0570 0.8920 ;
        RECT 0.7350 0.8920 2.0570 0.9420 ;
        RECT 1.6470 0.9420 1.6970 1.5640 ;
        RECT 1.9510 0.9420 2.0010 1.5650 ;
        RECT 0.7350 0.9420 0.7850 1.5640 ;
        RECT 1.0390 0.9420 1.0890 1.5640 ;
        RECT 1.3430 0.9420 1.3930 1.5640 ;
    END
    ANTENNADIFFAREA 0.6952 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 2.3950 1.7730 ;
    LAYER M1 ;
      RECT 0.6390 0.6600 1.9560 0.7100 ;
      RECT 0.2790 0.5020 0.3290 0.5370 ;
      RECT 0.2790 0.1160 0.3290 0.5760 ;
      RECT 0.2790 0.8920 0.3290 1.5640 ;
      RECT 0.2790 0.5370 0.6730 0.5870 ;
      RECT 0.3290 0.9310 0.6330 0.9390 ;
      RECT 0.5830 0.8920 0.6330 1.5640 ;
      RECT 0.2790 0.8920 0.6330 0.9310 ;
      RECT 0.5830 0.1160 0.6330 0.5760 ;
      RECT 0.3290 0.9390 0.5830 0.9420 ;
      RECT 0.6080 0.8920 0.6850 0.9420 ;
      RECT 0.6390 0.8420 0.6850 0.8500 ;
      RECT 0.6350 0.8500 0.6850 0.8920 ;
      RECT 0.6350 0.5370 0.6850 0.6100 ;
      RECT 0.6380 0.6100 0.6850 0.6370 ;
      RECT 0.6390 0.6420 0.6890 0.8420 ;
      RECT 0.6380 0.6370 0.6890 0.6420 ;
    LAYER PO ;
      RECT 0.0610 0.0710 0.0910 1.6060 ;
      RECT 0.5170 0.0690 0.5470 1.6060 ;
      RECT 1.8850 0.0690 1.9150 1.6060 ;
      RECT 2.0370 0.0690 2.0670 1.6060 ;
      RECT 2.1890 0.0690 2.2190 1.6060 ;
      RECT 0.2130 0.0710 0.2430 1.6060 ;
      RECT 0.3650 0.0690 0.3950 1.6060 ;
      RECT 1.7330 0.0690 1.7630 1.6060 ;
      RECT 1.5810 0.0690 1.6110 1.6060 ;
      RECT 1.4290 0.0690 1.4590 1.6060 ;
      RECT 0.6690 0.0690 0.6990 1.6060 ;
      RECT 0.8210 0.0690 0.8510 1.6060 ;
      RECT 1.2770 0.0690 1.3070 1.6060 ;
      RECT 1.1250 0.0690 1.1550 1.6060 ;
      RECT 0.9730 0.0690 1.0030 1.6060 ;
  END
END NBUFFX8_LVT

MACRO NMT1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.76 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.0970 0.3590 0.2070 ;
        RECT 0.2790 0.2070 0.3290 0.4750 ;
    END
    ANTENNADIFFAREA 0.0428 ;
    ANTENNAGATEAREA 0.0428 ;
  END S

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 0.7600 0.0300 ;
    END
  END VSS

  PIN D
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 0.4010 0.5110 0.5110 ;
        RECT 0.4310 0.1170 0.4810 0.4010 ;
    END
    ANTENNADIFFAREA 0.0428 ;
  END D

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.3590 0.5830 ;
        RECT 0.2490 0.5830 0.4210 0.6330 ;
        RECT 0.2490 0.6330 0.3590 0.6630 ;
    END
    ANTENNAGATEAREA 0.0126 ;
  END G

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 0.7600 1.7020 ;
    END
  END VDD
  OBS
    LAYER NWELL ;
      RECT -0.1250 0.6790 0.8650 1.7730 ;
    LAYER PO ;
      RECT 0.6690 0.0670 0.6990 0.6490 ;
      RECT 0.2130 0.0670 0.2430 0.6490 ;
      RECT 0.0610 0.0670 0.0910 0.6490 ;
      RECT 0.5170 0.0670 0.5470 0.6490 ;
      RECT 0.3650 0.0670 0.3950 0.6490 ;
  END
END NMT1_LVT

MACRO NMT2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.912 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5830 0.1510 0.6330 0.4010 ;
        RECT 0.5530 0.4010 0.6630 0.4600 ;
        RECT 0.2790 0.4600 0.6630 0.5100 ;
        RECT 0.2790 0.1510 0.3290 0.4600 ;
        RECT 0.5530 0.5100 0.6630 0.5110 ;
    END
    ANTENNADIFFAREA 0.0856 ;
    ANTENNAGATEAREA 0.0856 ;
  END S

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 0.9120 1.7020 ;
    END
  END VDD

  PIN D
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 0.0970 0.5110 0.2070 ;
        RECT 0.4310 0.2070 0.4810 0.3250 ;
    END
    ANTENNADIFFAREA 0.0512 ;
  END D

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 0.9120 0.0300 ;
    END
  END VSS

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 0.7050 0.5110 0.8150 ;
        RECT 0.4310 0.6400 0.4810 0.7050 ;
        RECT 0.3390 0.5900 0.5730 0.6400 ;
    END
    ANTENNAGATEAREA 0.0252 ;
  END G
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.0270 1.7730 ;
    LAYER PO ;
      RECT 0.5170 0.0740 0.5470 0.6560 ;
      RECT 0.3650 0.0740 0.3950 0.6560 ;
      RECT 0.6690 0.0740 0.6990 0.6560 ;
      RECT 0.0610 0.0740 0.0910 0.6560 ;
      RECT 0.2130 0.0780 0.2430 0.6560 ;
      RECT 0.8210 0.0740 0.8510 0.6560 ;
  END
END NMT2_LVT

MACRO NMT3_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.216 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.5900 0.8770 0.6400 ;
        RECT 0.7050 0.6400 0.8150 0.6630 ;
        RECT 0.7050 0.5530 0.8150 0.5900 ;
    END
    ANTENNAGATEAREA 0.0504 ;
  END G

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.2160 0.0300 ;
    END
  END VSS

  PIN D
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4310 0.1390 0.8150 0.1890 ;
        RECT 0.4310 0.1240 0.4810 0.1390 ;
        RECT 0.7050 0.0970 0.8150 0.1390 ;
        RECT 0.7050 0.1890 0.8150 0.2210 ;
        RECT 0.4310 0.1890 0.4810 0.3130 ;
        RECT 0.7350 0.2210 0.7850 0.3130 ;
    END
    ANTENNADIFFAREA 0.1024 ;
  END D

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.2160 1.7020 ;
    END
  END VDD

  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2790 0.1240 0.3290 0.4530 ;
        RECT 0.2790 0.4530 0.9670 0.5030 ;
        RECT 0.8570 0.4010 0.9670 0.4530 ;
        RECT 0.8570 0.5030 0.9670 0.5110 ;
        RECT 0.5830 0.3010 0.6330 0.4530 ;
        RECT 0.8870 0.1240 0.9370 0.4010 ;
    END
    ANTENNADIFFAREA 0.1368 ;
    ANTENNAGATEAREA 0.1368 ;
  END S
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.3310 1.7730 ;
    LAYER PO ;
      RECT 0.9730 0.0740 1.0030 0.6560 ;
      RECT 0.5170 0.0740 0.5470 0.6560 ;
      RECT 0.8210 0.0740 0.8510 0.6560 ;
      RECT 0.0610 0.0740 0.0910 0.6560 ;
      RECT 0.2130 0.0740 0.2430 0.6560 ;
      RECT 1.1250 0.0740 1.1550 0.6560 ;
      RECT 0.3650 0.0740 0.3950 0.6560 ;
      RECT 0.6690 0.0740 0.6990 0.6560 ;
  END
END NMT3_LVT

MACRO LSUPX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.128 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6200 2.2130 1.1810 2.2630 ;
        RECT 1.0090 2.2630 1.1190 2.3350 ;
    END
    ANTENNAGATEAREA 0.0444 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.2700 1.2710 1.2710 ;
        RECT 1.0390 1.2200 1.2710 1.2700 ;
        RECT 1.0390 1.2700 1.0890 1.5670 ;
        RECT 1.1210 1.1610 1.2710 1.2200 ;
        RECT 1.1210 1.0330 1.1710 1.1610 ;
        RECT 1.0390 0.9830 1.1710 1.0330 ;
        RECT 1.0390 0.1260 1.0890 0.9830 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.1280 1.7020 ;
        RECT 1.7700 1.7020 1.8800 1.7760 ;
        RECT 1.7700 1.5690 1.8800 1.6420 ;
        RECT 0.4310 1.3380 0.4810 1.6420 ;
        RECT 1.4950 1.3030 1.5450 1.6420 ;
        RECT 0.5820 1.3520 0.6320 1.6420 ;
        RECT 0.8870 1.2000 0.9370 1.6420 ;
        RECT 1.0390 1.7020 1.0890 2.0230 ;
    END
  END VSS

  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.1280 0.0300 ;
        RECT 0.8870 0.0300 0.9370 0.9440 ;
        RECT 1.4950 0.0300 1.5450 0.5260 ;
        RECT 0.4310 0.0300 0.4810 0.8240 ;
        RECT 0.5830 0.0300 0.6330 0.8240 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 2.1280 3.3740 ;
    END
  END VDDH

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 3.0100 2.1280 3.0700 ;
        RECT 1.3140 3.0700 1.4240 3.1440 ;
        RECT 1.3140 2.9370 1.4240 3.0100 ;
        RECT 1.0390 2.5350 1.0890 3.0100 ;
        RECT 1.3430 2.4280 1.3930 2.9370 ;
    END
  END VDDL
  OBS
    LAYER NWELL ;
      RECT -0.1150 -0.1150 2.2430 0.9930 ;
      RECT -0.1150 3.2240 2.2430 3.4590 ;
      RECT 2.0080 2.3510 2.2430 3.2240 ;
      RECT -0.1150 2.3510 0.1150 3.2240 ;
      RECT 0.5750 2.2320 1.4790 2.7640 ;
    LAYER M1 ;
      RECT 0.7340 1.0840 1.0310 1.1330 ;
      RECT 0.7660 1.0830 1.0310 1.0840 ;
      RECT 0.7750 0.9340 0.8250 1.0830 ;
      RECT 0.7340 1.1330 0.8250 1.1340 ;
      RECT 0.3390 0.8840 0.8250 0.9340 ;
      RECT 0.7350 1.1340 0.7850 1.5840 ;
      RECT 0.7350 0.5580 0.7850 0.8840 ;
      RECT 0.2390 0.9840 0.7250 1.0340 ;
      RECT 0.2800 1.0340 0.3300 1.5840 ;
      RECT 0.2390 0.8310 0.2890 0.9840 ;
      RECT 0.2390 0.7810 0.3290 0.8310 ;
      RECT 0.2790 0.5580 0.3290 0.7810 ;
      RECT 0.8870 2.4230 1.2810 2.4730 ;
      RECT 1.1910 2.4730 1.2410 2.7090 ;
      RECT 0.3330 2.1110 1.2810 2.1610 ;
      RECT 1.1920 1.9870 1.2420 2.1110 ;
      RECT 1.2310 2.1610 1.2810 2.4230 ;
      RECT 0.8870 2.4730 0.9370 2.7090 ;
      RECT 0.8870 1.9870 0.9370 2.1110 ;
    LAYER PO ;
      RECT 2.0370 0.0740 2.0670 2.7800 ;
      RECT 0.2130 0.0890 0.2430 2.7800 ;
      RECT 0.5170 0.0890 0.5470 2.7800 ;
      RECT 0.0610 0.0890 0.0910 2.7800 ;
      RECT 0.8210 0.0780 0.8510 2.7800 ;
      RECT 0.6690 1.1880 0.6990 2.7810 ;
      RECT 1.5810 0.0740 1.6110 2.7800 ;
      RECT 1.2770 0.0750 1.3070 2.7800 ;
      RECT 0.6690 0.0890 0.6990 1.0450 ;
      RECT 0.3650 0.0890 0.3950 0.9380 ;
      RECT 1.4290 0.0690 1.4590 2.7800 ;
      RECT 1.1250 0.0870 1.1550 2.7780 ;
      RECT 0.3650 1.1680 0.3950 2.7800 ;
      RECT 1.8850 0.0740 1.9150 2.7800 ;
      RECT 0.9730 0.0560 1.0030 1.7660 ;
      RECT 1.7330 0.0740 1.7630 2.7800 ;
      RECT 0.9730 1.8810 1.0030 2.7810 ;
  END
END LSUPX1_LVT

MACRO LSUPX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.28 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 3.0100 2.2800 3.0700 ;
        RECT 1.7700 3.0700 1.8800 3.1440 ;
        RECT 1.7700 2.9370 1.8800 3.0100 ;
        RECT 1.3430 2.4280 1.3930 3.0100 ;
        RECT 1.0390 2.5350 1.0890 3.0100 ;
    END
  END VDDL

  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.2800 0.0300 ;
        RECT 0.5830 0.0300 0.6330 0.4230 ;
        RECT 0.4310 0.0300 0.4810 0.7910 ;
        RECT 1.9510 0.0300 2.0010 0.5260 ;
        RECT 1.1910 0.0300 1.2410 0.9360 ;
        RECT 1.6470 0.0300 1.6970 0.8440 ;
        RECT 0.5830 0.4230 0.9370 0.4730 ;
        RECT 0.8870 0.4730 0.9370 0.8020 ;
        RECT 0.5830 0.4730 0.6330 0.7910 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 2.2800 3.3740 ;
    END
  END VDDH

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.2800 1.7020 ;
        RECT 1.9220 1.7020 2.0320 1.7760 ;
        RECT 1.9220 1.5690 2.0320 1.6420 ;
        RECT 1.0390 1.7020 1.0890 2.0230 ;
        RECT 0.8870 1.2600 0.9370 1.6420 ;
        RECT 1.6470 1.2780 1.6970 1.6420 ;
        RECT 0.5820 1.2600 0.6320 1.6420 ;
        RECT 0.4310 1.2460 0.4810 1.6420 ;
        RECT 1.1910 1.2980 1.2410 1.6420 ;
        RECT 1.9510 1.3030 2.0010 1.5690 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7990 1.1000 1.9940 1.1500 ;
        RECT 1.9440 0.9670 1.9940 1.1000 ;
        RECT 1.7990 1.1500 1.8490 1.1780 ;
        RECT 1.9200 0.9510 2.0310 0.9670 ;
        RECT 1.4940 1.1780 1.8490 1.2280 ;
        RECT 1.4950 0.9010 2.0310 0.9510 ;
        RECT 1.4950 1.2280 1.5450 1.5360 ;
        RECT 1.7990 1.2280 1.8490 1.5360 ;
        RECT 1.4950 0.1180 1.5450 0.9010 ;
        RECT 1.9200 0.8570 2.0310 0.9010 ;
        RECT 1.7990 0.1180 1.8490 0.9010 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6310 2.2130 1.1810 2.2630 ;
        RECT 1.0090 2.2630 1.1190 2.3350 ;
    END
    ANTENNAGATEAREA 0.0474 ;
  END A
  OBS
    LAYER NWELL ;
      RECT -0.1150 3.2240 2.3950 3.4590 ;
      RECT -0.1150 2.3510 0.1150 3.2240 ;
      RECT 2.1570 2.3510 2.3900 3.2240 ;
      RECT 0.5900 2.2340 1.4790 2.7640 ;
      RECT -0.1150 -0.1510 2.3950 0.9930 ;
    LAYER M1 ;
      RECT 0.7660 1.0830 1.0310 1.0840 ;
      RECT 0.7340 1.0840 1.0310 1.1330 ;
      RECT 0.7750 0.9010 0.8250 1.0830 ;
      RECT 0.7340 1.1330 0.8250 1.1340 ;
      RECT 0.3390 0.8510 0.8250 0.9010 ;
      RECT 0.7350 1.1340 0.7850 1.5130 ;
      RECT 0.7350 0.5250 0.7850 0.8510 ;
      RECT 1.0810 1.1820 1.3330 1.1830 ;
      RECT 1.0390 1.1830 1.3330 1.2320 ;
      RECT 1.0810 1.0330 1.1310 1.1820 ;
      RECT 1.0390 1.2320 1.1310 1.2330 ;
      RECT 1.0390 0.9830 1.1310 1.0330 ;
      RECT 1.0390 1.2330 1.0890 1.5670 ;
      RECT 1.0390 0.6280 1.0890 0.9830 ;
      RECT 0.3330 2.1110 1.2810 2.1610 ;
      RECT 1.1920 1.9870 1.2420 2.1110 ;
      RECT 1.1910 2.3620 1.2410 2.4230 ;
      RECT 0.8870 2.4230 1.2410 2.4730 ;
      RECT 1.1910 2.4730 1.2410 2.7090 ;
      RECT 1.1910 2.3130 1.2810 2.3620 ;
      RECT 1.2310 2.1610 1.2810 2.3130 ;
      RECT 0.8870 1.9870 0.9370 2.1110 ;
      RECT 0.8870 2.4730 0.9370 2.7090 ;
      RECT 0.2390 0.9840 0.7250 1.0340 ;
      RECT 0.2800 1.0340 0.3300 1.5760 ;
      RECT 0.2390 0.7980 0.2890 0.9840 ;
      RECT 0.2390 0.7480 0.3290 0.7980 ;
      RECT 0.2790 0.5250 0.3290 0.7480 ;
      RECT 1.3430 1.0010 1.7890 1.0370 ;
      RECT 1.3440 1.0370 1.7890 1.0500 ;
      RECT 1.3440 1.0500 1.7490 1.0510 ;
      RECT 1.3830 1.0510 1.4330 1.2810 ;
      RECT 1.3430 0.1180 1.3930 1.0010 ;
      RECT 1.3430 1.2810 1.4330 1.3310 ;
      RECT 1.3430 1.3310 1.3930 1.5640 ;
    LAYER PO ;
      RECT 0.0610 0.0890 0.0910 2.7800 ;
      RECT 0.5170 0.0890 0.5470 2.7800 ;
      RECT 0.2130 0.0890 0.2430 2.7800 ;
      RECT 0.9730 1.8810 1.0030 2.7810 ;
      RECT 0.9730 0.0790 1.0030 1.7660 ;
      RECT 2.1890 0.0740 2.2190 2.7800 ;
      RECT 0.3650 1.1680 0.3950 2.7800 ;
      RECT 1.1250 0.0870 1.1550 2.7780 ;
      RECT 1.8850 0.0690 1.9150 2.7800 ;
      RECT 1.7330 0.0620 1.7630 2.7730 ;
      RECT 0.3650 0.0900 0.3950 0.9050 ;
      RECT 0.6690 0.0890 0.6990 1.0450 ;
      RECT 1.4290 0.0690 1.4590 2.7800 ;
      RECT 1.2770 0.0680 1.3070 2.7730 ;
      RECT 2.0370 0.0740 2.0670 2.7800 ;
      RECT 1.5810 0.0620 1.6110 2.7730 ;
      RECT 0.6690 1.1880 0.6990 2.7810 ;
      RECT 0.8210 0.0780 0.8510 2.7800 ;
  END
END LSUPX2_LVT

MACRO LSUPX4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.584 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6310 2.2130 1.1810 2.2630 ;
        RECT 1.0090 2.2630 1.1190 2.3350 ;
    END
    ANTENNAGATEAREA 0.051 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4950 0.8940 2.3420 0.9440 ;
        RECT 1.4950 0.1180 1.5450 0.8940 ;
        RECT 2.1030 0.1180 2.1530 0.8940 ;
        RECT 1.7990 0.1180 1.8490 0.8940 ;
        RECT 2.2240 0.9440 2.3420 0.9670 ;
        RECT 2.2240 0.8570 2.3420 0.8940 ;
        RECT 2.2920 0.9670 2.3420 1.1410 ;
        RECT 2.2920 0.8550 2.3420 0.8570 ;
        RECT 1.4940 1.1410 2.3420 1.1910 ;
        RECT 2.1030 1.1910 2.1530 1.5360 ;
        RECT 1.7990 1.1910 1.8490 1.5360 ;
        RECT 1.4950 1.1910 1.5450 1.5360 ;
    END
    ANTENNADIFFAREA 0.3976 ;
  END Y

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.5840 1.7020 ;
        RECT 2.2260 1.7020 2.3360 1.7760 ;
        RECT 2.2260 1.5690 2.3360 1.6420 ;
        RECT 0.8870 1.2600 0.9370 1.6420 ;
        RECT 1.0390 1.7020 1.0890 2.0230 ;
        RECT 1.9510 1.2780 2.0010 1.6420 ;
        RECT 1.1910 1.2980 1.2410 1.6420 ;
        RECT 0.4310 1.1540 0.4810 1.6420 ;
        RECT 0.5820 1.1680 0.6320 1.6420 ;
        RECT 1.6470 1.2770 1.6970 1.6420 ;
        RECT 2.2550 1.3030 2.3050 1.5690 ;
    END
  END VSS

  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.5840 0.0300 ;
        RECT 1.9510 0.0300 2.0010 0.8440 ;
        RECT 1.6470 0.0300 1.6970 0.8440 ;
        RECT 1.1910 0.0300 1.2410 0.9360 ;
        RECT 0.8870 0.0300 0.9370 0.7190 ;
        RECT 2.2540 0.0300 2.3040 0.5260 ;
        RECT 0.4310 0.0300 0.4810 0.6780 ;
        RECT 0.5830 0.0300 0.6330 0.6780 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 2.5840 3.3740 ;
    END
  END VDDH

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 3.0100 2.5840 3.0700 ;
        RECT 1.6180 3.0700 1.7280 3.1440 ;
        RECT 1.6180 2.9370 1.7280 3.0100 ;
        RECT 1.0390 2.5350 1.0890 3.0100 ;
        RECT 1.3430 2.4280 1.3930 3.0100 ;
    END
  END VDDL
  OBS
    LAYER NWELL ;
      RECT -0.1150 -0.1150 2.6990 0.9930 ;
      RECT -0.1150 3.2240 2.6990 3.4590 ;
      RECT 2.4690 2.3510 2.6990 3.2240 ;
      RECT -0.1150 2.3510 0.1150 3.2240 ;
      RECT 0.5750 2.2340 1.4800 2.7640 ;
    LAYER M1 ;
      RECT 1.3430 2.1610 1.3930 2.3180 ;
      RECT 1.1910 2.3180 1.3930 2.3680 ;
      RECT 0.3330 2.1110 1.3930 2.1610 ;
      RECT 0.8870 1.9870 0.9370 2.1110 ;
      RECT 0.8870 2.4730 0.9370 2.7090 ;
      RECT 1.1910 2.3680 1.2410 2.4230 ;
      RECT 1.1920 1.9870 1.2420 2.1110 ;
      RECT 0.8870 2.4230 1.2410 2.4730 ;
      RECT 1.1910 2.4730 1.2410 2.7090 ;
      RECT 0.7660 1.0830 1.0290 1.0840 ;
      RECT 0.7340 1.0840 1.0290 1.1330 ;
      RECT 0.7750 0.7880 0.8250 1.0830 ;
      RECT 0.7340 1.1330 0.8250 1.1340 ;
      RECT 0.3390 0.7380 0.8250 0.7880 ;
      RECT 0.7350 1.1340 0.7850 1.5680 ;
      RECT 0.7350 0.4120 0.7850 0.7380 ;
      RECT 1.0810 1.1820 1.3330 1.1830 ;
      RECT 1.0390 1.1830 1.3330 1.2320 ;
      RECT 1.0810 1.0330 1.1310 1.1820 ;
      RECT 1.0390 1.2320 1.1310 1.2330 ;
      RECT 1.0390 0.9830 1.1310 1.0330 ;
      RECT 1.0390 1.2330 1.0890 1.5560 ;
      RECT 1.0390 0.5480 1.0890 0.9830 ;
      RECT 1.3430 1.0010 2.0930 1.0510 ;
      RECT 1.3430 0.1180 1.3930 1.0010 ;
      RECT 1.3830 1.0510 1.4330 1.2810 ;
      RECT 1.3430 1.2810 1.4330 1.3310 ;
      RECT 1.3430 1.3310 1.3930 1.5640 ;
      RECT 0.2390 0.8380 0.7250 0.8880 ;
      RECT 0.2800 0.8880 0.3300 1.5680 ;
      RECT 0.2390 0.6850 0.2890 0.8380 ;
      RECT 0.2390 0.6350 0.3290 0.6850 ;
      RECT 0.2790 0.4120 0.3290 0.6350 ;
    LAYER PO ;
      RECT 1.8850 0.0680 1.9150 2.7800 ;
      RECT 2.0370 0.0680 2.0670 2.7800 ;
      RECT 0.2130 0.0890 0.2430 2.7800 ;
      RECT 0.5170 0.0890 0.5470 2.7800 ;
      RECT 0.0610 0.0890 0.0910 2.7800 ;
      RECT 0.8210 0.0780 0.8510 2.7800 ;
      RECT 0.6690 1.0680 0.6990 2.7810 ;
      RECT 1.5810 0.0680 1.6110 2.7800 ;
      RECT 2.3410 0.0740 2.3710 2.7800 ;
      RECT 1.2770 0.0680 1.3070 2.7800 ;
      RECT 1.4290 0.0680 1.4590 2.7800 ;
      RECT 0.6690 0.0910 0.6990 0.9280 ;
      RECT 0.3650 0.0880 0.3950 0.9010 ;
      RECT 1.7330 0.0680 1.7630 2.7800 ;
      RECT 2.1890 0.0680 2.2190 2.7800 ;
      RECT 1.1250 0.0870 1.1550 2.7780 ;
      RECT 0.3650 1.0680 0.3950 2.7800 ;
      RECT 2.4930 0.0740 2.5230 2.7800 ;
      RECT 0.9730 0.0790 1.0030 1.7660 ;
      RECT 0.9730 1.8810 1.0030 2.7810 ;
  END
END LSUPX4_LVT

MACRO LSUPX8_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.344 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6310 2.2130 1.1810 2.2630 ;
        RECT 1.0090 2.2630 1.1190 2.3350 ;
    END
    ANTENNAGATEAREA 0.051 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6470 1.1330 2.9850 1.1830 ;
        RECT 1.9510 1.1830 2.0010 1.5360 ;
        RECT 1.6470 1.1830 1.6970 1.5360 ;
        RECT 2.2550 1.1830 2.3050 1.5360 ;
        RECT 2.8630 1.1830 2.9130 1.5360 ;
        RECT 2.5590 1.1830 2.6090 1.5360 ;
        RECT 2.9350 0.9680 2.9850 1.1330 ;
        RECT 2.9350 0.9440 3.0950 0.9680 ;
        RECT 1.6480 0.9190 3.0950 0.9440 ;
        RECT 1.6470 0.8940 3.0950 0.9190 ;
        RECT 2.9850 0.8570 3.0950 0.8940 ;
        RECT 2.8630 0.1180 2.9130 0.8940 ;
        RECT 2.5590 0.1180 2.6090 0.8940 ;
        RECT 2.2550 0.1180 2.3050 0.8940 ;
        RECT 1.9510 0.1180 2.0010 0.8940 ;
        RECT 1.6470 0.1180 1.6970 0.8940 ;
    END
    ANTENNADIFFAREA 0.6952 ;
  END Y

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.3440 1.7020 ;
        RECT 2.9860 1.7020 3.0960 1.7760 ;
        RECT 2.9860 1.5690 3.0960 1.6420 ;
        RECT 1.4950 1.2980 1.5450 1.6420 ;
        RECT 1.1910 1.2980 1.2410 1.6420 ;
        RECT 0.4310 1.1440 0.4810 1.6420 ;
        RECT 0.8870 1.2000 0.9370 1.6420 ;
        RECT 0.5820 1.1570 0.6320 1.6420 ;
        RECT 2.1030 1.2790 2.1530 1.6420 ;
        RECT 2.4070 1.2790 2.4570 1.6420 ;
        RECT 1.7990 1.2780 1.8490 1.6420 ;
        RECT 2.7110 1.2990 2.7610 1.6420 ;
        RECT 1.0390 1.7020 1.0890 1.9950 ;
        RECT 3.0150 1.3030 3.0650 1.5690 ;
    END
  END VSS

  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.3440 0.0300 ;
        RECT 2.4070 0.0300 2.4570 0.8440 ;
        RECT 1.7990 0.0300 1.8490 0.8440 ;
        RECT 0.8870 0.0300 0.9370 0.7370 ;
        RECT 2.1030 0.0300 2.1530 0.8440 ;
        RECT 2.7110 0.0300 2.7610 0.8440 ;
        RECT 1.1910 0.0300 1.2410 0.9360 ;
        RECT 3.0150 0.0300 3.0650 0.5260 ;
        RECT 0.4310 0.0300 0.4810 0.6820 ;
        RECT 0.5830 0.0300 0.6330 0.6820 ;
        RECT 1.4950 0.0300 1.5450 0.9360 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 3.3440 3.3740 ;
    END
  END VDDH

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 3.0100 3.3440 3.0700 ;
        RECT 2.2260 3.0700 2.3360 3.1440 ;
        RECT 2.2260 2.9370 2.3360 3.0100 ;
        RECT 1.0390 2.5350 1.0890 3.0100 ;
        RECT 1.3430 2.4280 1.3930 3.0100 ;
    END
  END VDDL
  OBS
    LAYER NWELL ;
      RECT -0.1150 -0.1150 3.4590 0.9930 ;
      RECT -0.1150 3.2240 3.4590 3.4590 ;
      RECT 3.2290 2.3510 3.4590 3.2240 ;
      RECT -0.1150 2.3510 0.1150 3.2240 ;
      RECT 0.5750 2.2340 1.6170 2.7640 ;
    LAYER M1 ;
      RECT 0.7350 1.0840 1.0290 1.1340 ;
      RECT 0.7350 1.1340 0.7850 1.5830 ;
      RECT 0.7750 0.7920 0.8250 1.0840 ;
      RECT 0.3390 0.7420 0.8250 0.7920 ;
      RECT 0.7350 0.4160 0.7850 0.7420 ;
      RECT 1.0390 1.1860 1.3330 1.2360 ;
      RECT 1.0390 1.2360 1.0890 1.5480 ;
      RECT 1.0390 1.1850 1.1290 1.1860 ;
      RECT 1.0790 1.0340 1.1290 1.1850 ;
      RECT 1.0390 0.9830 1.1290 1.0340 ;
      RECT 1.0390 0.5650 1.0890 0.9830 ;
      RECT 0.2390 0.8420 0.7250 0.8920 ;
      RECT 0.2800 0.8920 0.3300 1.5840 ;
      RECT 0.2390 0.6890 0.2890 0.8420 ;
      RECT 0.2390 0.6390 0.3290 0.6890 ;
      RECT 0.2790 0.4160 0.3290 0.6390 ;
      RECT 0.3330 2.0830 1.2810 2.1330 ;
      RECT 1.1920 1.9590 1.2420 2.0830 ;
      RECT 1.1910 2.4350 1.2410 2.7090 ;
      RECT 1.2310 2.1330 1.2810 2.3850 ;
      RECT 0.8870 2.3850 1.2810 2.4350 ;
      RECT 0.8870 1.9590 0.9370 2.0830 ;
      RECT 0.8870 2.4350 0.9370 2.7090 ;
      RECT 1.3430 1.0330 2.8530 1.0830 ;
      RECT 1.3430 0.1180 1.3930 1.0330 ;
      RECT 1.3830 1.0830 1.4330 1.2870 ;
      RECT 1.3430 1.2870 1.4330 1.3370 ;
      RECT 1.3430 1.3370 1.3930 1.5640 ;
      RECT 1.2510 1.7810 1.4850 1.8310 ;
    LAYER PO ;
      RECT 0.6690 1.0570 0.6990 2.7810 ;
      RECT 1.7330 0.0680 1.7630 2.7800 ;
      RECT 3.1010 0.0740 3.1310 2.7800 ;
      RECT 1.4290 0.0680 1.4590 2.7800 ;
      RECT 1.2770 0.0680 1.3070 2.7800 ;
      RECT 1.5810 0.0690 1.6110 2.7800 ;
      RECT 0.3650 0.1150 0.3950 0.9130 ;
      RECT 1.8850 0.0680 1.9150 2.7800 ;
      RECT 0.9730 0.0790 1.0030 1.7380 ;
      RECT 2.9490 0.0690 2.9790 2.7800 ;
      RECT 1.1250 0.0870 1.1550 2.7780 ;
      RECT 0.3650 1.0580 0.3950 2.7800 ;
      RECT 2.7970 0.0680 2.8270 2.7800 ;
      RECT 2.6450 0.0680 2.6750 2.7800 ;
      RECT 2.4930 0.0680 2.5230 2.7800 ;
      RECT 2.3410 0.0680 2.3710 2.7800 ;
      RECT 2.1890 0.0680 2.2190 2.7800 ;
      RECT 2.0370 0.0680 2.0670 2.7800 ;
      RECT 0.9730 1.8530 1.0030 2.7810 ;
      RECT 3.2530 0.0740 3.2830 2.7800 ;
      RECT 0.6690 0.1020 0.6990 0.9030 ;
      RECT 0.2130 0.1140 0.2430 2.7800 ;
      RECT 0.5170 0.0890 0.5470 2.7800 ;
      RECT 0.0610 0.1140 0.0910 2.7800 ;
      RECT 0.8210 0.0780 0.8510 2.7800 ;
  END
END LSUPX8_LVT

MACRO MUX21X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.976 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.9760 0.0300 ;
        RECT 1.4950 0.0300 1.5450 0.5580 ;
        RECT 0.5830 0.0300 0.6330 0.2950 ;
        RECT 0.8870 0.0300 0.9370 0.2960 ;
        RECT 1.0390 0.0300 1.0890 0.2960 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.9760 1.7020 ;
        RECT 0.8870 1.3850 0.9370 1.6420 ;
        RECT 1.0390 1.3850 1.0890 1.6420 ;
        RECT 1.4950 1.3850 1.5450 1.6420 ;
        RECT 0.5830 1.3850 0.6330 1.6420 ;
    END
  END VDD

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.4150 0.6630 ;
        RECT 0.3550 0.6630 0.4050 0.6920 ;
        RECT 0.3550 0.4990 0.4050 0.5530 ;
    END
    ANTENNAGATEAREA 0.0189 ;
  END A1

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5070 0.7290 0.9670 0.7790 ;
        RECT 0.8110 0.7790 0.9670 0.8150 ;
        RECT 0.8110 0.7050 0.9670 0.7290 ;
        RECT 0.5070 0.7790 0.5570 1.1540 ;
        RECT 0.9170 0.6640 0.9670 0.7050 ;
        RECT 0.9170 0.6140 1.1650 0.6640 ;
        RECT 1.1150 0.6640 1.1650 0.6960 ;
    END
    ANTENNAGATEAREA 0.0378 ;
  END S0

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6470 0.1520 1.6970 0.5080 ;
        RECT 1.6470 0.5080 1.8010 0.5580 ;
        RECT 1.7510 0.5580 1.8010 0.7050 ;
        RECT 1.7510 0.7050 1.8800 0.7650 ;
        RECT 1.6470 0.7650 1.8800 0.8150 ;
        RECT 1.6470 0.8150 1.6970 1.5500 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2510 1.0090 1.4230 1.1190 ;
    END
    ANTENNAGATEAREA 0.0189 ;
  END A2
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 2.0910 1.7730 ;
    LAYER M1 ;
      RECT 1.1150 0.7520 1.2930 0.8020 ;
      RECT 1.2430 0.5640 1.2930 0.7520 ;
      RECT 0.5070 0.5140 1.2930 0.5640 ;
      RECT 1.1150 0.8020 1.1650 1.0740 ;
      RECT 0.7350 1.0740 1.1650 1.1240 ;
      RECT 0.5070 0.4240 0.5570 0.5140 ;
      RECT 0.7350 0.1610 0.7850 0.5140 ;
      RECT 0.7350 1.1240 0.7850 1.2320 ;
      RECT 1.3430 0.6080 1.6520 0.6580 ;
      RECT 1.5140 0.6580 1.5640 1.2850 ;
      RECT 0.2790 1.2850 1.5640 1.3350 ;
      RECT 1.3430 0.1390 1.3930 0.6080 ;
      RECT 1.3430 1.3350 1.3930 1.5500 ;
      RECT 0.2790 1.3350 0.3290 1.5490 ;
      RECT 0.2790 0.9440 0.3290 1.2850 ;
      RECT 0.1490 0.8940 0.3290 0.9440 ;
      RECT 0.1490 0.2870 0.3290 0.3370 ;
      RECT 0.2790 0.1380 0.3290 0.2870 ;
      RECT 0.1490 0.3370 0.1990 0.8940 ;
    LAYER PO ;
      RECT 1.1250 0.0720 1.1550 0.7110 ;
      RECT 0.0610 0.0710 0.0910 1.6090 ;
      RECT 0.3650 0.0690 0.3950 1.6090 ;
      RECT 0.2130 0.0710 0.2430 1.6090 ;
      RECT 1.5810 0.0720 1.6110 1.6100 ;
      RECT 1.7330 0.0720 1.7630 1.6100 ;
      RECT 1.8850 0.0720 1.9150 1.6100 ;
      RECT 0.6690 0.0710 0.6990 1.6090 ;
      RECT 0.5170 0.0710 0.5470 0.5250 ;
      RECT 0.8210 0.0720 0.8510 1.6100 ;
      RECT 1.1250 1.0150 1.1550 1.6100 ;
      RECT 0.9730 0.0720 1.0030 1.6100 ;
      RECT 1.2770 0.0720 1.3070 1.6100 ;
      RECT 1.4290 0.0720 1.4590 1.6100 ;
      RECT 0.5170 1.0050 0.5470 1.6090 ;
  END
END MUX21X1_LVT

MACRO MUX21X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.128 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.1280 0.0300 ;
        RECT 1.7990 0.0300 1.8490 0.3290 ;
        RECT 1.4950 0.0300 1.5450 0.4980 ;
        RECT 1.0390 0.0300 1.0890 0.3880 ;
        RECT 0.8870 0.0300 0.9370 0.3880 ;
        RECT 0.5830 0.0300 0.6330 0.3870 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6470 0.1320 1.6970 0.4480 ;
        RECT 1.6470 0.4480 1.9480 0.4980 ;
        RECT 1.8980 0.4980 1.9480 0.7050 ;
        RECT 1.8980 0.7050 2.0310 0.8150 ;
        RECT 1.8980 0.8150 1.9480 0.8350 ;
        RECT 1.6470 0.8350 1.9480 0.8850 ;
        RECT 1.6470 0.8850 1.6970 1.5450 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.1280 1.7020 ;
        RECT 1.4950 1.2790 1.5450 1.6420 ;
        RECT 1.7990 1.0030 1.8490 1.6420 ;
        RECT 0.5830 1.2920 0.6330 1.6420 ;
        RECT 1.0390 1.2730 1.0890 1.6420 ;
        RECT 0.8870 1.2920 0.9370 1.6420 ;
    END
  END VDD

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5070 0.7050 0.9670 0.7550 ;
        RECT 0.5070 0.6630 0.5570 0.7050 ;
        RECT 0.8110 0.7550 0.9670 0.8150 ;
        RECT 0.9170 0.6640 0.9670 0.7050 ;
        RECT 0.5070 0.7550 0.5570 1.0290 ;
        RECT 0.9170 0.6140 1.1650 0.6640 ;
        RECT 1.1150 0.6640 1.1650 0.6960 ;
    END
    ANTENNAGATEAREA 0.0468 ;
  END S0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2300 0.5530 0.4150 0.6630 ;
        RECT 0.3550 0.6630 0.4050 0.6920 ;
        RECT 0.3550 0.4990 0.4050 0.5530 ;
    END
    ANTENNAGATEAREA 0.0234 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2510 0.8570 1.4230 0.9670 ;
    END
    ANTENNAGATEAREA 0.0234 ;
  END A2
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 2.2430 1.7730 ;
    LAYER M1 ;
      RECT 1.2430 0.5640 1.2930 0.7460 ;
      RECT 0.5070 0.5140 1.2930 0.5640 ;
      RECT 1.1150 0.7460 1.2930 0.7960 ;
      RECT 1.1150 0.7960 1.1650 0.9800 ;
      RECT 0.7350 0.9800 1.1650 1.0060 ;
      RECT 0.7350 1.0060 1.1640 1.0300 ;
      RECT 0.5070 0.5090 0.5570 0.5140 ;
      RECT 0.5070 0.5640 0.5570 0.6130 ;
      RECT 0.7350 0.1440 0.7850 0.5140 ;
      RECT 0.7350 1.0300 0.7850 1.1220 ;
      RECT 1.3430 0.6100 1.7890 0.6600 ;
      RECT 1.3430 0.1240 1.3930 0.6100 ;
      RECT 1.3430 1.2220 1.3930 1.5500 ;
      RECT 1.5380 0.6600 1.5880 1.1720 ;
      RECT 0.2790 1.1720 1.5880 1.2220 ;
      RECT 0.2790 1.2220 0.3290 1.5490 ;
      RECT 0.2790 0.9440 0.3290 1.1720 ;
      RECT 0.0970 0.8940 0.3290 0.9440 ;
      RECT 0.0970 0.3740 0.3290 0.4240 ;
      RECT 0.2790 0.1380 0.3290 0.3740 ;
      RECT 0.0970 0.4240 0.1470 0.8940 ;
    LAYER PO ;
      RECT 1.1250 0.0720 1.1550 0.7110 ;
      RECT 2.0370 0.0580 2.0670 1.5960 ;
      RECT 1.8850 0.0580 1.9150 1.5960 ;
      RECT 1.7330 0.0720 1.7630 1.6040 ;
      RECT 1.5810 0.0720 1.6110 1.6100 ;
      RECT 0.5170 0.8950 0.5470 1.6090 ;
      RECT 1.4290 0.0720 1.4590 1.6100 ;
      RECT 1.2770 0.0720 1.3070 1.6100 ;
      RECT 0.9730 0.0720 1.0030 1.6100 ;
      RECT 1.1250 0.8930 1.1550 1.6100 ;
      RECT 0.8210 0.0720 0.8510 1.6100 ;
      RECT 0.5170 0.0710 0.5470 0.6270 ;
      RECT 0.6690 0.0710 0.6990 1.6090 ;
      RECT 0.2130 0.0710 0.2430 1.6090 ;
      RECT 0.3650 0.0690 0.3950 1.6090 ;
      RECT 0.0610 0.0710 0.0910 1.6090 ;
  END
END MUX21X2_LVT

MACRO MUX41X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.344 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.1400 0.6660 3.2480 0.8420 ;
        RECT 3.1400 0.4530 3.1900 0.6660 ;
        RECT 3.1400 0.8420 3.1900 0.9210 ;
        RECT 3.0150 0.4030 3.1900 0.4530 ;
        RECT 3.0150 0.9210 3.1900 0.9710 ;
        RECT 3.0150 0.2160 3.0650 0.4030 ;
        RECT 3.0150 0.9710 3.0650 1.1460 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7070 0.0970 1.8790 0.2070 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END A1

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.1620 1.4440 2.7080 1.4940 ;
        RECT 2.5290 1.4940 2.6590 1.5810 ;
    END
    ANTENNAGATEAREA 0.048 ;
  END S0

  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6590 0.2720 1.1400 0.3220 ;
        RECT 0.6590 0.1300 0.7090 0.2720 ;
        RECT 1.0900 0.1300 1.1400 0.2720 ;
        RECT 0.2490 0.0800 0.7250 0.1300 ;
        RECT 1.0900 0.0800 1.4850 0.1300 ;
        RECT 0.2490 0.1300 0.4170 0.2070 ;
    END
    ANTENNAGATEAREA 0.072 ;
  END S1

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 0.8210 1.0370 0.8710 ;
        RECT 0.8570 0.8710 0.9670 0.9670 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END A3

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7950 0.5530 0.9670 0.6690 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END A4

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4650 0.7050 1.6370 0.8280 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END A2

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.3440 0.0300 ;
        RECT 0.1310 0.0300 0.1810 0.4120 ;
        RECT 1.5350 0.0300 1.5850 0.2570 ;
        RECT 2.8630 0.0300 2.9130 0.2210 ;
        RECT 0.9280 0.0300 0.9780 0.1720 ;
        RECT 2.7600 0.0300 2.8100 0.1920 ;
        RECT 0.1310 0.4120 0.3290 0.4620 ;
        RECT 1.5350 0.2570 1.7130 0.3070 ;
        RECT 0.8670 0.1720 0.9780 0.2220 ;
        RECT 2.5430 0.1920 2.8100 0.2420 ;
        RECT 0.2790 0.4620 0.3290 0.6250 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.3440 1.7020 ;
        RECT 0.2790 1.0500 0.3290 1.6420 ;
        RECT 0.8870 1.3350 0.9370 1.6420 ;
        RECT 1.6470 1.3200 1.6970 1.6420 ;
        RECT 3.0970 1.4880 3.1470 1.6420 ;
        RECT 2.8630 1.4380 3.1470 1.4880 ;
        RECT 2.8630 1.2580 2.9130 1.4380 ;
        RECT 2.5430 1.2080 2.9130 1.2580 ;
    END
  END VDD
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 3.4590 1.7730 ;
    LAYER M1 ;
      RECT 1.4430 1.1200 1.7530 1.1700 ;
      RECT 1.7030 0.7560 1.7530 1.1200 ;
      RECT 1.7030 0.7060 1.9060 0.7560 ;
      RECT 1.8560 0.7000 1.9060 0.7060 ;
      RECT 1.8560 0.6500 1.9410 0.7000 ;
      RECT 0.6830 1.1850 0.7330 1.4420 ;
      RECT 0.4310 1.4420 0.7330 1.4920 ;
      RECT 0.4310 0.4720 0.4810 1.4420 ;
      RECT 1.4430 1.1700 1.4930 1.3760 ;
      RECT 1.1150 1.3760 1.4930 1.4260 ;
      RECT 1.4010 1.4260 1.4930 1.4780 ;
      RECT 1.1150 1.1850 1.1650 1.3760 ;
      RECT 0.6830 1.1350 1.1650 1.1850 ;
      RECT 1.0690 0.9720 1.1190 1.1350 ;
      RECT 1.0690 0.9220 1.1650 0.9720 ;
      RECT 1.1150 0.5490 1.1650 0.9220 ;
      RECT 1.9350 0.9110 2.0450 0.9610 ;
      RECT 1.9950 0.5080 2.0450 0.9110 ;
      RECT 1.3430 0.4580 2.1530 0.5080 ;
      RECT 2.1030 0.5080 2.1530 0.8800 ;
      RECT 1.3430 0.5080 1.3930 1.3100 ;
      RECT 2.4010 1.1040 2.7610 1.1540 ;
      RECT 2.7110 0.3920 2.7610 1.1040 ;
      RECT 2.4010 1.1540 2.4510 1.3440 ;
      RECT 2.0560 1.3440 2.4510 1.3940 ;
      RECT 2.0560 1.3940 2.1060 1.4280 ;
      RECT 2.0090 1.4280 2.1060 1.4780 ;
      RECT 2.8780 0.6580 3.0050 0.7080 ;
      RECT 2.2550 0.9330 2.6340 0.9830 ;
      RECT 2.5840 0.3420 2.6340 0.9330 ;
      RECT 2.2550 0.4920 2.3050 0.9330 ;
      RECT 2.5840 0.2920 2.9280 0.3420 ;
      RECT 2.8780 0.3420 2.9280 0.6580 ;
      RECT 1.1150 1.5260 1.1650 1.5780 ;
      RECT 0.9870 1.4760 1.1650 1.5260 ;
      RECT 0.9870 1.2850 1.0370 1.4760 ;
      RECT 0.7830 1.2350 1.0370 1.2850 ;
      RECT 0.7830 1.2850 0.8330 1.5420 ;
      RECT 0.4850 1.5420 0.8330 1.5920 ;
      RECT 2.4070 0.4070 2.4570 0.8800 ;
      RECT 0.5830 0.3840 2.4570 0.4070 ;
      RECT 1.2190 0.3570 2.4570 0.3840 ;
      RECT 0.5830 0.4340 0.6330 1.3920 ;
      RECT 0.5830 0.4070 1.2690 0.4340 ;
      RECT 1.2190 0.4340 1.2690 1.0350 ;
      RECT 1.1690 1.0350 1.2690 1.0850 ;
      RECT 1.8030 0.8560 1.8530 1.2200 ;
      RECT 1.8030 0.8060 1.9410 0.8560 ;
      RECT 1.5470 1.2200 1.8530 1.2700 ;
      RECT 1.5470 1.2700 1.5970 1.5420 ;
      RECT 1.2450 1.5420 1.5970 1.5920 ;
      RECT 2.0040 0.0800 2.2450 0.1300 ;
      RECT 2.3150 0.0800 2.7010 0.1300 ;
    LAYER PO ;
      RECT 1.7330 0.0710 1.7630 1.6090 ;
      RECT 2.1890 0.7480 2.2190 1.6090 ;
      RECT 2.1890 0.0690 2.2190 0.6480 ;
      RECT 1.4290 0.0710 1.4590 0.6730 ;
      RECT 1.4290 0.8320 1.4590 1.6090 ;
      RECT 0.5170 0.0710 0.5470 1.6090 ;
      RECT 0.2130 0.0710 0.2430 1.6090 ;
      RECT 3.1010 0.0720 3.1310 1.6100 ;
      RECT 0.9730 0.0710 1.0030 1.6090 ;
      RECT 2.6450 0.0720 2.6750 1.6100 ;
      RECT 1.8850 0.0710 1.9150 0.7000 ;
      RECT 1.8850 0.8070 1.9150 1.6090 ;
      RECT 2.3410 0.0690 2.3710 0.6240 ;
      RECT 2.7970 0.0720 2.8270 1.6100 ;
      RECT 1.1250 0.0710 1.1550 0.6270 ;
      RECT 1.2770 0.0720 1.3070 1.6100 ;
      RECT 1.1250 0.7560 1.1550 1.6090 ;
      RECT 0.6690 0.0710 0.6990 0.6270 ;
      RECT 3.2530 0.0720 3.2830 1.6100 ;
      RECT 0.0610 0.0710 0.0910 1.6090 ;
      RECT 2.0370 0.0690 2.0670 1.6090 ;
      RECT 0.6690 0.7500 0.6990 1.6090 ;
      RECT 0.3650 0.0710 0.3950 1.6090 ;
      RECT 2.9490 0.0720 2.9790 1.6100 ;
      RECT 2.3410 0.7480 2.3710 1.6090 ;
      RECT 0.8210 0.0710 0.8510 1.6090 ;
      RECT 2.4930 0.0710 2.5230 1.6090 ;
      RECT 1.5810 0.0710 1.6110 1.6090 ;
  END
END MUX41X1_LVT

MACRO MUX41X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.648 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2070 0.3660 3.2570 0.9210 ;
        RECT 2.9150 0.3160 3.2570 0.3660 ;
        RECT 2.8630 0.9210 3.2570 0.9710 ;
        RECT 2.9150 0.2850 2.9650 0.3160 ;
        RECT 3.1370 0.2490 3.2570 0.3160 ;
        RECT 3.1670 0.9710 3.2170 1.1460 ;
        RECT 2.8630 0.9710 2.9130 1.1460 ;
        RECT 2.8630 0.2350 2.9650 0.2850 ;
        RECT 2.8630 0.1790 2.9130 0.2350 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7110 0.0880 1.8560 0.2120 ;
    END
    ANTENNAGATEAREA 0.0264 ;
  END A1

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.1620 1.4440 2.7080 1.4940 ;
        RECT 2.5290 1.4940 2.6390 1.5750 ;
    END
    ANTENNAGATEAREA 0.0528 ;
  END S0

  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6590 0.2960 1.1400 0.3460 ;
        RECT 0.6590 0.1380 0.7090 0.2960 ;
        RECT 1.0900 0.1380 1.1400 0.2960 ;
        RECT 0.2490 0.0880 0.7250 0.1380 ;
        RECT 1.0900 0.0880 1.4850 0.1380 ;
        RECT 0.2490 0.1380 0.4170 0.2170 ;
    END
    ANTENNAGATEAREA 0.0792 ;
  END S1

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8490 0.8570 1.0250 0.9620 ;
        RECT 0.9630 0.7790 1.0130 0.8570 ;
    END
    ANTENNAGATEAREA 0.0264 ;
  END A3

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6930 0.5570 0.8690 0.7110 ;
    END
    ANTENNAGATEAREA 0.0264 ;
  END A4

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.6480 1.7020 ;
        RECT 0.2790 1.0500 0.3290 1.6420 ;
        RECT 0.8870 1.3270 0.9370 1.6420 ;
        RECT 1.6470 1.3100 1.6970 1.6420 ;
        RECT 3.0970 1.4880 3.1470 1.6420 ;
        RECT 2.8630 1.4380 3.1470 1.4880 ;
        RECT 2.8630 1.2580 2.9130 1.4380 ;
        RECT 2.5430 1.2080 2.9130 1.2580 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.6480 0.0300 ;
        RECT 0.1310 0.0300 0.1810 0.4120 ;
        RECT 1.5350 0.0300 1.5850 0.2620 ;
        RECT 3.0150 0.0300 3.0650 0.2660 ;
        RECT 0.8870 0.0300 0.9370 0.2460 ;
        RECT 2.7600 0.0300 2.8100 0.1940 ;
        RECT 0.1310 0.4120 0.3290 0.4620 ;
        RECT 1.5350 0.2620 1.7330 0.3120 ;
        RECT 2.5430 0.1940 2.8100 0.2440 ;
        RECT 0.2790 0.4620 0.3290 0.6250 ;
    END
  END VSS

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4650 0.7050 1.6370 0.8150 ;
    END
    ANTENNAGATEAREA 0.0264 ;
  END A2
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 3.7630 1.7730 ;
    LAYER M1 ;
      RECT 1.4430 1.1100 1.7530 1.1600 ;
      RECT 1.7030 0.6990 1.7530 1.1100 ;
      RECT 1.7030 0.6490 1.9410 0.6990 ;
      RECT 1.4430 1.1600 1.4930 1.3760 ;
      RECT 1.1150 1.3760 1.4930 1.4260 ;
      RECT 1.4190 1.4260 1.4690 1.4840 ;
      RECT 0.6830 1.1720 0.7330 1.4340 ;
      RECT 0.4310 1.4340 0.7330 1.4840 ;
      RECT 0.4310 0.4720 0.4810 1.4340 ;
      RECT 1.1150 1.1770 1.1650 1.3760 ;
      RECT 1.0750 1.1720 1.1650 1.1770 ;
      RECT 0.6830 1.1420 1.1650 1.1720 ;
      RECT 0.6840 1.1270 1.1650 1.1420 ;
      RECT 0.6840 1.1220 1.1250 1.1270 ;
      RECT 1.1150 0.5460 1.1650 0.9270 ;
      RECT 1.0500 0.4960 1.1650 0.5460 ;
      RECT 1.0750 0.9770 1.1250 1.1220 ;
      RECT 1.0750 0.9270 1.1650 0.9770 ;
      RECT 1.9350 0.9010 2.0450 0.9510 ;
      RECT 1.9950 0.5120 2.0450 0.9010 ;
      RECT 1.3430 0.4620 2.1530 0.5120 ;
      RECT 2.1030 0.5120 2.1530 0.8800 ;
      RECT 1.3430 0.5120 1.3930 1.3000 ;
      RECT 2.4010 1.1040 2.7610 1.1540 ;
      RECT 2.7110 0.4820 2.7610 1.1040 ;
      RECT 2.4010 1.1540 2.4510 1.3440 ;
      RECT 2.0560 1.3440 2.4510 1.3940 ;
      RECT 2.0560 1.3940 2.1060 1.4280 ;
      RECT 2.0090 1.4280 2.1060 1.4780 ;
      RECT 2.8110 0.6580 3.1570 0.7080 ;
      RECT 2.5840 0.4320 2.6340 0.9330 ;
      RECT 2.2550 0.9330 2.6340 0.9830 ;
      RECT 2.2550 0.4920 2.3050 0.9330 ;
      RECT 2.8110 0.4320 2.8610 0.6580 ;
      RECT 2.5840 0.3820 2.8610 0.4320 ;
      RECT 1.1150 1.5260 1.1650 1.5780 ;
      RECT 0.9870 1.4760 1.1650 1.5260 ;
      RECT 0.9870 1.2770 1.0370 1.4760 ;
      RECT 0.7830 1.2270 1.0370 1.2770 ;
      RECT 0.7830 1.2770 0.8330 1.5340 ;
      RECT 0.4850 1.5340 0.8330 1.5840 ;
      RECT 2.4070 0.4120 2.4570 0.8800 ;
      RECT 1.2190 0.3620 2.4570 0.3960 ;
      RECT 0.5830 0.3960 2.4570 0.4120 ;
      RECT 0.5830 0.4460 0.6330 1.3840 ;
      RECT 0.5830 0.4120 1.2690 0.4460 ;
      RECT 1.2190 0.4460 1.2690 1.0270 ;
      RECT 1.1750 1.0270 1.2690 1.0770 ;
      RECT 1.8030 0.8460 1.8530 1.2100 ;
      RECT 1.8030 0.7960 1.9410 0.8460 ;
      RECT 1.5470 1.2100 1.8530 1.2600 ;
      RECT 1.5470 1.2600 1.5970 1.5340 ;
      RECT 1.2450 1.5340 1.5970 1.5840 ;
      RECT 2.0040 0.0880 2.2450 0.1380 ;
      RECT 2.3150 0.0880 2.7010 0.1380 ;
    LAYER PO ;
      RECT 2.3410 0.7480 2.3710 1.6090 ;
      RECT 0.8210 0.0710 0.8510 1.6090 ;
      RECT 2.4930 0.0710 2.5230 1.6090 ;
      RECT 1.5810 0.0710 1.6110 1.6090 ;
      RECT 1.7330 0.0710 1.7630 1.6090 ;
      RECT 2.1890 0.7480 2.2190 1.6090 ;
      RECT 2.1890 0.0690 2.2190 0.6480 ;
      RECT 1.4290 0.0710 1.4590 0.6730 ;
      RECT 1.4290 0.8220 1.4590 1.6090 ;
      RECT 0.5170 0.0710 0.5470 1.6090 ;
      RECT 0.2130 0.0710 0.2430 1.6090 ;
      RECT 3.4050 0.0720 3.4350 1.6100 ;
      RECT 0.9730 0.0710 1.0030 1.6090 ;
      RECT 2.6450 0.0720 2.6750 1.6100 ;
      RECT 1.8850 0.0710 1.9150 0.6960 ;
      RECT 1.8850 0.7970 1.9150 1.6090 ;
      RECT 2.3410 0.0690 2.3710 0.6240 ;
      RECT 2.7970 0.0720 2.8270 1.6100 ;
      RECT 1.1250 0.0710 1.1550 0.6380 ;
      RECT 1.2770 0.0720 1.3070 1.6100 ;
      RECT 1.1250 0.7560 1.1550 1.6090 ;
      RECT 0.6690 0.0710 0.6990 0.6270 ;
      RECT 3.1010 0.0720 3.1310 1.6100 ;
      RECT 3.2530 0.0720 3.2830 1.6100 ;
      RECT 3.5570 0.0720 3.5870 1.6100 ;
      RECT 0.0610 0.0710 0.0910 1.6090 ;
      RECT 2.0370 0.0690 2.0670 1.6090 ;
      RECT 0.6690 0.7500 0.6990 1.6090 ;
      RECT 0.3650 0.0710 0.3950 1.6090 ;
      RECT 2.9490 0.0720 2.9790 1.6100 ;
  END
END MUX41X2_LVT

MACRO NAND2X0_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.912 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2540 0.7350 0.4260 0.7850 ;
        RECT 0.2540 0.7050 0.3590 0.7350 ;
        RECT 0.2540 0.7850 0.3590 0.8150 ;
    END
    ANTENNAGATEAREA 0.0186 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 1.0390 0.5730 1.0890 ;
        RECT 0.4010 1.0090 0.5060 1.0390 ;
        RECT 0.4010 1.0890 0.5060 1.1190 ;
    END
    ANTENNAGATEAREA 0.0186 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 0.8570 0.6730 0.9670 ;
        RECT 0.6230 0.9670 0.6730 1.1850 ;
        RECT 0.6230 0.6710 0.6730 0.8570 ;
        RECT 0.2790 1.1850 0.6730 1.2350 ;
        RECT 0.5830 0.6210 0.6730 0.6710 ;
        RECT 0.5830 1.2350 0.6330 1.5510 ;
        RECT 0.2790 1.2350 0.3290 1.5510 ;
        RECT 0.5830 0.1060 0.6330 0.6210 ;
    END
    ANTENNADIFFAREA 0.0938 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 0.9120 1.7020 ;
        RECT 0.4310 1.2850 0.4810 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 0.9120 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.4020 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.0270 1.7730 ;
    LAYER PO ;
      RECT 0.6690 0.0710 0.6990 1.6010 ;
      RECT 0.3650 0.0710 0.3950 1.6010 ;
      RECT 0.5170 0.0710 0.5470 1.6010 ;
      RECT 0.2130 0.0710 0.2430 1.6010 ;
      RECT 0.8210 0.0710 0.8510 1.6010 ;
      RECT 0.0610 0.0710 0.0910 1.6010 ;
  END
END NAND2X0_LVT

MACRO NAND2X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.52 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4560 0.8870 0.6630 0.9370 ;
        RECT 0.5530 0.9370 0.6630 0.9670 ;
        RECT 0.5530 0.8570 0.6630 0.8870 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6880 0.4250 0.8180 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END A2

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 0.8540 1.2810 0.9670 ;
        RECT 1.1910 0.9670 1.2410 1.5610 ;
        RECT 1.2310 0.5250 1.2810 0.8540 ;
        RECT 1.1910 0.4750 1.2810 0.5250 ;
        RECT 1.1910 0.1340 1.2410 0.4750 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0280 1.5200 0.0280 ;
        RECT 0.2790 0.0280 0.3290 0.4790 ;
        RECT 1.0390 0.0280 1.0890 0.3160 ;
        RECT 0.7350 0.0280 0.7850 0.3110 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6440 1.5200 1.7000 ;
        RECT 0.4310 1.1930 0.4810 1.6440 ;
        RECT 1.0390 1.1880 1.0890 1.6440 ;
        RECT 0.7350 1.1830 0.7850 1.6440 ;
    END
  END VDD
  OBS
    LAYER NWELL ;
      RECT -0.0910 0.6790 1.6110 1.7810 ;
    LAYER M1 ;
      RECT 0.9270 0.6420 1.1810 0.6920 ;
      RECT 0.9270 0.6920 0.9770 0.8560 ;
      RECT 0.9270 0.5050 0.9770 0.6420 ;
      RECT 0.8870 0.8560 0.9770 0.9060 ;
      RECT 0.8870 0.4550 0.9770 0.5050 ;
      RECT 0.8870 0.9060 0.9370 1.5560 ;
      RECT 0.8870 0.1290 0.9370 0.4550 ;
      RECT 0.7130 0.7310 0.8770 0.7810 ;
      RECT 0.7130 0.6630 0.7630 0.7310 ;
      RECT 0.5830 0.6130 0.7630 0.6630 ;
      RECT 0.7130 0.7810 0.7630 1.0830 ;
      RECT 0.2790 1.0830 0.7630 1.1330 ;
      RECT 0.2790 1.1330 0.3290 1.5510 ;
      RECT 0.5830 1.1330 0.6330 1.5510 ;
      RECT 0.5830 0.1060 0.6330 0.6130 ;
    LAYER PO ;
      RECT 1.1250 0.0640 1.1550 1.6070 ;
      RECT 0.8210 0.0640 0.8510 1.6020 ;
      RECT 1.4290 0.0640 1.4590 1.6000 ;
      RECT 1.2770 0.0640 1.3070 1.6050 ;
      RECT 0.9730 0.0640 1.0030 1.6050 ;
      RECT 0.0610 0.0710 0.0910 1.6010 ;
      RECT 0.2130 0.0710 0.2430 1.6010 ;
      RECT 0.5170 0.0710 0.5470 1.6010 ;
      RECT 0.3650 0.0710 0.3950 1.6010 ;
      RECT 0.6690 0.0710 0.6990 1.6010 ;
  END
END NAND2X1_LVT

MACRO NAND2X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.672 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.7350 0.5110 0.7850 ;
        RECT 0.4010 0.7850 0.5110 0.8150 ;
        RECT 0.4010 0.7050 0.5110 0.7350 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END A2

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.6720 0.0300 ;
        RECT 0.7350 0.0300 0.7850 0.3150 ;
        RECT 1.0390 0.0300 1.0890 0.4860 ;
        RECT 1.3430 0.0300 1.3930 0.4860 ;
        RECT 0.2790 0.0300 0.3290 0.4790 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1910 0.5530 1.5750 0.5920 ;
        RECT 1.4650 0.5920 1.5750 0.6630 ;
        RECT 1.1910 0.5420 1.5150 0.5530 ;
        RECT 1.4650 0.6630 1.5150 0.7420 ;
        RECT 1.1910 0.1200 1.2410 0.5420 ;
        RECT 1.1910 0.7420 1.5150 0.7920 ;
        RECT 1.1910 0.7920 1.2410 1.5560 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.6720 1.7020 ;
        RECT 0.7350 1.1830 0.7850 1.6420 ;
        RECT 1.0390 0.8150 1.0890 1.6420 ;
        RECT 1.3430 0.9070 1.3930 1.6420 ;
        RECT 0.4310 1.1930 0.4810 1.6420 ;
    END
  END VDD

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4560 0.8870 0.6630 0.9370 ;
        RECT 0.5530 0.9370 0.6630 0.9670 ;
        RECT 0.5530 0.8570 0.6630 0.8870 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END A1
  OBS
    LAYER NWELL ;
      RECT -0.0910 0.6790 1.7630 1.7730 ;
    LAYER M1 ;
      RECT 0.7100 0.7310 0.8770 0.7810 ;
      RECT 0.7130 0.6630 0.7630 0.7310 ;
      RECT 0.5830 0.6130 0.7630 0.6630 ;
      RECT 0.2790 1.0830 0.7630 1.1330 ;
      RECT 0.5830 0.1210 0.6330 0.6130 ;
      RECT 0.5830 1.1330 0.6330 1.5510 ;
      RECT 0.7130 0.7810 0.7630 1.0830 ;
      RECT 0.2790 1.1330 0.3290 1.5510 ;
      RECT 0.9270 0.6420 1.3330 0.6920 ;
      RECT 0.9270 0.6920 0.9770 0.8560 ;
      RECT 0.9270 0.5050 0.9770 0.6420 ;
      RECT 0.8870 0.8560 0.9770 0.9060 ;
      RECT 0.8870 0.4550 0.9770 0.5050 ;
      RECT 0.8870 0.9060 0.9370 1.5560 ;
      RECT 0.8870 0.1330 0.9370 0.4550 ;
    LAYER PO ;
      RECT 0.6690 0.0710 0.6990 1.6010 ;
      RECT 0.3650 0.0710 0.3950 1.6010 ;
      RECT 0.5170 0.0710 0.5470 1.6010 ;
      RECT 0.2130 0.0710 0.2430 1.6010 ;
      RECT 0.0610 0.0710 0.0910 1.6010 ;
      RECT 1.2770 0.0640 1.3070 1.6070 ;
      RECT 0.9730 0.0640 1.0030 1.6000 ;
      RECT 0.8210 0.0640 0.8510 1.6100 ;
      RECT 1.1250 0.0640 1.1550 1.6080 ;
      RECT 1.5810 0.0640 1.6110 1.6000 ;
      RECT 1.4290 0.0640 1.4590 1.6020 ;
  END
END NAND2X2_LVT

MACRO NAND2X4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.976 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.7350 0.5110 0.7850 ;
        RECT 0.4010 0.7850 0.5110 0.8150 ;
        RECT 0.4010 0.7050 0.5110 0.7350 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END A2

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.9760 0.0300 ;
        RECT 0.7350 0.0300 0.7850 0.5170 ;
        RECT 1.1910 0.0300 1.2410 0.3970 ;
        RECT 1.4950 0.0300 1.5450 0.3970 ;
        RECT 0.2790 0.0300 0.3290 0.4870 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0390 0.1310 1.0890 0.5130 ;
        RECT 1.0390 0.5130 1.8020 0.5530 ;
        RECT 1.3430 0.1310 1.3930 0.5130 ;
        RECT 1.6470 0.1310 1.6970 0.5130 ;
        RECT 1.0390 0.5530 1.8890 0.5630 ;
        RECT 1.7520 0.5630 1.8890 0.6630 ;
        RECT 1.7520 0.6630 1.8020 0.7430 ;
        RECT 1.0390 0.7430 1.8020 0.7930 ;
        RECT 1.0390 0.7930 1.0890 1.5650 ;
        RECT 1.3430 0.7930 1.3930 1.5650 ;
        RECT 1.6470 0.7930 1.6970 1.5650 ;
    END
    ANTENNADIFFAREA 0.3972 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.9760 1.7020 ;
        RECT 0.7350 0.8230 0.7850 1.6420 ;
        RECT 0.4310 1.2470 0.4810 1.6420 ;
        RECT 1.1910 0.9160 1.2410 1.6420 ;
        RECT 1.4950 0.9160 1.5450 1.6420 ;
    END
  END VDD

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4910 0.8870 0.6630 0.9370 ;
        RECT 0.5530 0.9370 0.6630 0.9670 ;
        RECT 0.5530 0.8570 0.6630 0.8870 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END A1
  OBS
    LAYER NWELL ;
      RECT -0.0910 0.6790 2.0690 1.7810 ;
    LAYER M1 ;
      RECT 0.9270 0.6420 1.6370 0.6920 ;
      RECT 0.9270 0.5370 0.9770 0.6420 ;
      RECT 0.9270 0.6920 0.9770 0.7080 ;
      RECT 0.8870 0.4870 0.9770 0.5370 ;
      RECT 0.8870 0.7080 0.9770 0.7580 ;
      RECT 0.8870 0.1310 0.9370 0.4870 ;
      RECT 0.8870 0.7580 0.9370 1.5640 ;
      RECT 0.2380 0.6050 0.8770 0.6550 ;
      RECT 0.5830 0.1310 0.6330 0.6050 ;
      RECT 0.2380 1.1010 0.6330 1.1510 ;
      RECT 0.5830 1.1510 0.6330 1.5590 ;
      RECT 0.2380 0.6550 0.2880 1.1010 ;
      RECT 0.2790 1.1510 0.3290 1.5590 ;
    LAYER PO ;
      RECT 0.6690 0.0710 0.6990 1.6010 ;
      RECT 0.3650 0.0710 0.3950 1.6090 ;
      RECT 0.5170 0.0710 0.5470 1.6090 ;
      RECT 0.2130 0.0710 0.2430 1.6090 ;
      RECT 0.0610 0.0710 0.0910 1.6010 ;
      RECT 1.2770 0.0710 1.3070 1.6100 ;
      RECT 1.4290 0.0710 1.4590 1.6100 ;
      RECT 1.5810 0.0710 1.6110 1.6100 ;
      RECT 1.8850 0.0720 1.9150 1.6100 ;
      RECT 1.7330 0.0720 1.7630 1.6100 ;
      RECT 1.1250 0.0710 1.1550 1.6100 ;
      RECT 0.9730 0.0640 1.0030 1.6080 ;
      RECT 0.8210 0.0640 0.8510 1.6100 ;
  END
END NAND2X4_LVT

MACRO NAND3X0_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.064 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8550 0.8570 0.9650 0.9670 ;
        RECT 0.8650 0.6550 0.9150 0.8570 ;
        RECT 0.8650 0.9670 0.9150 1.0900 ;
        RECT 0.7350 0.6050 0.9150 0.6550 ;
        RECT 0.4560 1.0900 0.9150 1.0910 ;
        RECT 0.7350 0.1060 0.7850 0.6050 ;
        RECT 0.4310 1.0910 0.9150 1.1400 ;
        RECT 0.4310 1.1400 0.4810 1.5510 ;
        RECT 0.7350 1.1400 0.7850 1.5510 ;
    END
    ANTENNADIFFAREA 0.1348 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6430 0.7350 0.8150 0.7850 ;
        RECT 0.7050 0.7850 0.8150 0.8150 ;
        RECT 0.7050 0.7050 0.8150 0.7350 ;
    END
    ANTENNAGATEAREA 0.0246 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4910 0.8870 0.6630 0.9370 ;
        RECT 0.5530 0.9370 0.6630 0.9670 ;
        RECT 0.5530 0.8570 0.6630 0.8870 ;
    END
    ANTENNAGATEAREA 0.0246 ;
  END A2

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.0640 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.4790 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.0640 1.7020 ;
        RECT 0.2790 1.1930 0.3290 1.6420 ;
        RECT 0.5830 1.1930 0.6330 1.6420 ;
    END
  END VDD

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.8570 0.3590 0.8870 ;
        RECT 0.2490 0.8870 0.4210 0.9370 ;
        RECT 0.2490 0.9370 0.3590 0.9670 ;
    END
    ANTENNAGATEAREA 0.0246 ;
  END A3
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.1780 1.7730 ;
    LAYER PO ;
      RECT 0.0610 0.0710 0.0910 1.6100 ;
      RECT 0.8210 0.0710 0.8510 1.6100 ;
      RECT 0.2130 0.0710 0.2430 1.6100 ;
      RECT 0.5170 0.0710 0.5470 1.6100 ;
      RECT 0.3650 0.0710 0.3950 1.6100 ;
      RECT 0.6690 0.0710 0.6990 1.6100 ;
      RECT 0.9730 0.0710 1.0030 1.6100 ;
  END
END NAND3X0_LVT

MACRO LSDNSSX8_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.584 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.5840 0.0300 ;
        RECT 0.7350 0.0300 0.7850 0.4100 ;
        RECT 1.7990 0.0300 1.8490 0.4100 ;
        RECT 2.1030 0.0300 2.1530 0.4100 ;
        RECT 1.4950 0.0300 1.5450 0.4100 ;
        RECT 0.4310 0.0300 0.4810 0.4100 ;
        RECT 1.1910 0.0300 1.2410 0.4100 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6600 0.8770 0.7100 ;
        RECT 0.2490 0.7100 0.3620 0.8150 ;
    END
    ANTENNAGATEAREA 0.0312 ;
  END A

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.5840 1.7020 ;
        RECT 0.7350 0.9920 0.7850 1.6420 ;
        RECT 1.7990 0.9920 1.8490 1.6420 ;
        RECT 2.1030 0.9920 2.1530 1.6420 ;
        RECT 1.4950 0.9920 1.5450 1.6420 ;
        RECT 1.1910 0.9920 1.2410 1.6420 ;
        RECT 0.4310 0.9920 0.4810 1.6420 ;
    END
  END VDDL

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0390 0.5370 2.4870 0.5870 ;
        RECT 2.3110 0.5870 2.4870 0.6630 ;
        RECT 1.9510 0.3150 2.0010 0.5370 ;
        RECT 2.2550 0.3160 2.3050 0.5370 ;
        RECT 1.6470 0.3150 1.6970 0.5370 ;
        RECT 1.0390 0.3150 1.0890 0.5370 ;
        RECT 1.3430 0.3150 1.3930 0.5370 ;
        RECT 2.3110 0.6630 2.3610 0.8920 ;
        RECT 1.0390 0.8920 2.3610 0.9420 ;
        RECT 1.9510 0.9420 2.0010 1.5640 ;
        RECT 2.2550 0.9420 2.3050 1.5650 ;
        RECT 1.0390 0.9420 1.0890 1.5640 ;
        RECT 1.3430 0.9420 1.3930 1.5640 ;
        RECT 1.6470 0.9420 1.6970 1.5640 ;
    END
    ANTENNADIFFAREA 0.6044 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 2.6990 1.7730 ;
    LAYER M1 ;
      RECT 0.9270 0.6600 2.2600 0.7100 ;
      RECT 0.2790 0.8920 0.3290 1.5640 ;
      RECT 0.2790 0.5020 0.3290 0.5370 ;
      RECT 0.2790 0.3150 0.3290 0.5760 ;
      RECT 0.5830 0.8920 0.6330 1.5640 ;
      RECT 0.5830 0.3150 0.6330 0.5760 ;
      RECT 0.2790 0.8920 0.9370 0.9310 ;
      RECT 0.9120 0.8920 0.9770 0.9420 ;
      RECT 0.8870 0.8920 0.9370 1.5640 ;
      RECT 0.8870 0.3150 0.9370 0.5760 ;
      RECT 0.2790 0.5370 0.9650 0.5870 ;
      RECT 0.9270 0.5370 0.9770 0.9420 ;
      RECT 0.3290 0.9310 0.9370 0.9420 ;
    LAYER PO ;
      RECT 0.3650 0.0710 0.3950 1.6060 ;
      RECT 0.8210 0.0690 0.8510 1.6060 ;
      RECT 0.2130 0.0710 0.2430 1.6060 ;
      RECT 2.1890 0.0690 2.2190 1.6060 ;
      RECT 2.3410 0.0690 2.3710 1.6060 ;
      RECT 2.4930 0.0690 2.5230 1.6060 ;
      RECT 0.5170 0.0710 0.5470 1.6060 ;
      RECT 0.6690 0.0690 0.6990 1.6060 ;
      RECT 2.0370 0.0690 2.0670 1.6060 ;
      RECT 1.8850 0.0690 1.9150 1.6060 ;
      RECT 1.7330 0.0690 1.7630 1.6060 ;
      RECT 0.0610 0.0710 0.0910 1.6060 ;
      RECT 0.9730 0.0690 1.0030 1.6060 ;
      RECT 1.1250 0.0690 1.1550 1.6060 ;
      RECT 1.5810 0.0690 1.6110 1.6060 ;
      RECT 1.4290 0.0690 1.4590 1.6060 ;
      RECT 1.2770 0.0690 1.3070 1.6060 ;
  END
END LSDNSSX8_LVT

MACRO LSDNX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.128 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 3.0100 2.1280 3.0700 ;
        RECT 0.8580 3.0700 0.9680 3.1430 ;
        RECT 0.8580 2.9360 0.9680 3.0100 ;
        RECT 1.1910 2.5200 1.2410 3.0100 ;
        RECT 0.8830 2.3430 0.9390 2.9360 ;
    END
  END VDDH

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.1280 0.0300 ;
        RECT 0.2760 0.0300 0.3320 0.7690 ;
        RECT 0.5800 0.0300 0.6360 0.7520 ;
        RECT 1.1880 0.0300 1.2440 0.5040 ;
        RECT 0.8840 0.0300 0.9400 0.8370 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 2.1280 3.3740 ;
    END
  END VDDL

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.1280 1.7020 ;
        RECT 0.2760 1.3050 0.3320 1.6420 ;
        RECT 1.6180 1.7020 1.7280 1.7750 ;
        RECT 1.6180 1.5680 1.7280 1.6420 ;
        RECT 1.1880 1.2700 1.2440 1.6420 ;
        RECT 0.5800 1.1880 0.6360 1.6420 ;
        RECT 0.8840 1.1700 0.9400 1.6420 ;
        RECT 0.8840 1.7020 0.9400 2.0070 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0370 1.0760 1.1830 1.1320 ;
        RECT 1.1270 0.8680 1.1830 1.0760 ;
        RECT 1.0370 1.1320 1.0930 1.5700 ;
        RECT 1.1270 0.8670 1.3100 0.8680 ;
        RECT 1.0360 0.8110 1.3100 0.8670 ;
        RECT 1.0360 0.1880 1.0920 0.8110 ;
        RECT 1.1610 0.7050 1.3100 0.8110 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7940 2.2070 1.1410 2.2630 ;
        RECT 0.9970 2.2630 1.1410 2.3370 ;
        RECT 0.9970 2.2030 1.1410 2.2070 ;
    END
    ANTENNAGATEAREA 0.0132 ;
  END A
  OBS
    LAYER NWELL ;
      RECT -0.1150 3.2240 2.2430 3.4590 ;
      RECT -0.1150 2.3510 0.1150 3.2240 ;
      RECT 2.0130 2.3510 2.2430 3.2240 ;
      RECT 0.5750 2.2340 1.4250 2.7640 ;
      RECT -0.1150 -0.1150 2.2430 0.9930 ;
    LAYER M1 ;
      RECT 0.7750 0.9670 1.0290 1.0230 ;
      RECT 0.7750 1.0230 0.8310 1.0810 ;
      RECT 0.7750 0.9140 0.8310 0.9670 ;
      RECT 0.7320 1.0810 0.8310 1.1370 ;
      RECT 0.7330 0.8580 0.8310 0.9140 ;
      RECT 0.7320 1.1370 0.7880 1.4860 ;
      RECT 0.7330 0.1310 0.7890 0.8580 ;
      RECT 0.4820 0.9670 0.7250 1.0230 ;
      RECT 0.4820 1.0230 0.5380 1.0910 ;
      RECT 0.4820 0.9090 0.5380 0.9670 ;
      RECT 0.4200 0.8530 0.5380 0.9090 ;
      RECT 0.4280 1.0910 0.5380 1.1380 ;
      RECT 0.4280 1.1380 0.5300 1.1470 ;
      RECT 0.4280 1.1470 0.4840 1.4430 ;
      RECT 0.4280 0.5070 0.4840 0.8530 ;
      RECT 0.1860 0.9670 0.4210 1.0230 ;
      RECT 0.7310 2.3710 0.7870 2.6410 ;
      RECT 0.6390 2.3150 0.7870 2.3710 ;
      RECT 0.6390 2.0790 0.7880 2.1350 ;
      RECT 0.7320 1.8600 0.7880 2.0790 ;
      RECT 0.6390 2.2620 0.6950 2.3150 ;
      RECT 0.3390 2.2060 0.6950 2.2620 ;
      RECT 0.6390 2.1350 0.6950 2.2060 ;
    LAYER PO ;
      RECT 1.7330 0.0690 1.7630 2.7800 ;
      RECT 0.3650 0.0890 0.3950 2.7800 ;
      RECT 1.1250 0.0870 1.1550 2.7780 ;
      RECT 1.8850 0.0690 1.9150 2.7800 ;
      RECT 1.5810 0.0690 1.6110 2.7800 ;
      RECT 1.2770 0.0750 1.3070 2.7800 ;
      RECT 1.4290 0.0750 1.4590 2.7800 ;
      RECT 2.0370 0.0740 2.0670 2.7800 ;
      RECT 0.9730 0.0680 1.0030 2.7800 ;
      RECT 0.8210 0.0780 0.8510 2.7800 ;
      RECT 0.0610 0.0890 0.0910 2.7800 ;
      RECT 0.6690 0.0890 0.6990 2.7810 ;
      RECT 0.5170 0.0890 0.5470 2.7800 ;
      RECT 0.2130 0.0890 0.2430 2.7800 ;
  END
END LSDNX1_LVT

MACRO LSDNX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.128 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 3.0100 2.1280 3.0700 ;
        RECT 1.6180 3.0700 1.7280 3.1430 ;
        RECT 1.6180 2.9360 1.7280 3.0100 ;
        RECT 0.8830 2.3430 0.9390 3.0100 ;
        RECT 1.1910 2.5200 1.2410 3.0100 ;
    END
  END VDDH

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.1280 0.0300 ;
        RECT 0.2760 0.0300 0.3320 0.8500 ;
        RECT 0.5800 0.0300 0.6360 0.7860 ;
        RECT 1.3400 0.0300 1.3960 0.4720 ;
        RECT 0.8870 0.0300 0.9370 0.7840 ;
        RECT 1.1890 0.0300 1.2450 0.7830 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 2.1280 3.3740 ;
    END
  END VDDL

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.1280 1.7020 ;
        RECT 0.2760 1.3050 0.3320 1.6420 ;
        RECT 1.6180 1.7020 1.7280 1.7750 ;
        RECT 1.6180 1.5680 1.7280 1.6420 ;
        RECT 0.5800 1.1880 0.6360 1.6420 ;
        RECT 1.3390 1.2680 1.3950 1.6420 ;
        RECT 1.1880 1.2020 1.2440 1.6420 ;
        RECT 0.8840 1.7020 0.9400 2.0250 ;
        RECT 0.8840 1.1540 0.9400 1.6420 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0360 1.0870 1.3370 1.1430 ;
        RECT 1.0360 1.1430 1.0920 1.5610 ;
        RECT 1.2810 0.9670 1.3370 1.0870 ;
        RECT 1.2810 0.9160 1.4780 0.9670 ;
        RECT 1.0360 0.8600 1.4780 0.9160 ;
        RECT 1.0360 0.1620 1.0920 0.8600 ;
        RECT 1.3130 0.7780 1.4780 0.8600 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7940 2.2070 1.1390 2.2630 ;
        RECT 0.9950 2.2630 1.1390 2.3350 ;
        RECT 0.9950 2.2010 1.1390 2.2070 ;
    END
    ANTENNAGATEAREA 0.0132 ;
  END A
  OBS
    LAYER NWELL ;
      RECT -0.1150 3.2240 2.2430 3.4590 ;
      RECT -0.1150 2.3510 0.1150 3.2240 ;
      RECT 2.0130 2.3510 2.2430 3.2240 ;
      RECT -0.1150 -0.1150 2.2430 1.0530 ;
      RECT 0.5750 2.2340 1.4250 2.7640 ;
    LAYER M1 ;
      RECT 0.7750 0.9790 1.1810 1.0350 ;
      RECT 0.7750 1.0350 0.8310 1.0810 ;
      RECT 0.7750 0.9140 0.8310 0.9790 ;
      RECT 0.7390 1.0810 0.8310 1.0820 ;
      RECT 0.7330 0.8580 0.8310 0.9140 ;
      RECT 0.7350 1.0820 0.8310 1.1370 ;
      RECT 0.7330 0.1310 0.7890 0.8580 ;
      RECT 0.7350 1.1370 0.7910 1.5620 ;
      RECT 0.4820 0.9670 0.7250 1.0230 ;
      RECT 0.4820 1.0230 0.5380 1.0910 ;
      RECT 0.4820 0.9090 0.5380 0.9670 ;
      RECT 0.4280 0.8530 0.5380 0.9090 ;
      RECT 0.4300 1.0910 0.5380 1.1380 ;
      RECT 0.4300 1.1380 0.5300 1.1470 ;
      RECT 0.4300 1.1470 0.4860 1.4430 ;
      RECT 0.4280 0.4260 0.4840 0.8530 ;
      RECT 0.1860 0.9670 0.4210 1.0230 ;
      RECT 0.7310 2.3710 0.7870 2.6410 ;
      RECT 0.6390 2.3150 0.7870 2.3710 ;
      RECT 0.6390 2.0790 0.7880 2.1350 ;
      RECT 0.7320 1.8810 0.7880 2.0790 ;
      RECT 0.6390 2.2620 0.6950 2.3150 ;
      RECT 0.3390 2.2060 0.6950 2.2620 ;
      RECT 0.6390 2.1350 0.6950 2.2060 ;
    LAYER PO ;
      RECT 1.7330 0.0690 1.7630 2.7800 ;
      RECT 0.3650 0.0890 0.3950 2.7800 ;
      RECT 1.1250 0.0530 1.1550 2.7780 ;
      RECT 1.8850 0.0690 1.9150 2.7800 ;
      RECT 1.5810 0.0690 1.6110 2.7800 ;
      RECT 1.2770 0.0750 1.3070 2.7800 ;
      RECT 1.4290 0.0750 1.4590 2.7800 ;
      RECT 2.0370 0.0740 2.0670 2.7800 ;
      RECT 0.9730 0.0530 1.0030 2.7800 ;
      RECT 0.8210 0.0780 0.8510 2.7800 ;
      RECT 0.0610 0.0890 0.0910 2.7800 ;
      RECT 0.6690 0.0890 0.6990 2.7810 ;
      RECT 0.5170 0.0890 0.5470 2.7800 ;
      RECT 0.2130 0.0890 0.2430 2.7800 ;
  END
END LSDNX2_LVT

MACRO LSDNX4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.128 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 3.0100 2.1280 3.0700 ;
        RECT 1.4660 3.0700 1.5760 3.1430 ;
        RECT 1.4660 2.9360 1.5760 3.0100 ;
        RECT 0.8830 2.3430 0.9390 3.0100 ;
        RECT 1.1910 2.5200 1.2410 3.0100 ;
    END
  END VDDH

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.1280 0.0300 ;
        RECT 0.2760 0.0300 0.3320 0.7880 ;
        RECT 1.0360 0.0300 1.0920 0.7450 ;
        RECT 1.3410 0.0300 1.3970 0.7450 ;
        RECT 0.5800 0.0300 0.6360 0.6730 ;
        RECT 1.6440 0.0300 1.7000 0.4820 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 2.1280 3.3740 ;
    END
  END VDDL

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.1280 1.7020 ;
        RECT 0.2500 1.7020 0.3600 1.7750 ;
        RECT 0.2500 1.5680 0.3600 1.6420 ;
        RECT 1.0360 1.2650 1.0920 1.6420 ;
        RECT 1.3400 1.2650 1.3960 1.6420 ;
        RECT 1.6440 1.2670 1.7000 1.6420 ;
        RECT 0.5800 1.1880 0.6360 1.6420 ;
        RECT 0.8840 1.7020 0.9400 2.0250 ;
        RECT 0.2760 1.3050 0.3320 1.5680 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8830 0.1050 0.9390 0.8460 ;
        RECT 0.8830 0.8460 1.7770 0.9020 ;
        RECT 1.6170 0.7780 1.7770 0.8460 ;
        RECT 1.4920 0.1570 1.5480 0.8460 ;
        RECT 1.1890 0.1570 1.2450 0.8460 ;
        RECT 1.5930 0.9020 1.7770 0.9670 ;
        RECT 1.5930 0.9670 1.6490 1.0850 ;
        RECT 0.8840 1.0850 1.6490 1.1410 ;
        RECT 0.8840 1.1410 0.9400 1.5530 ;
        RECT 1.4920 1.1410 1.5480 1.5560 ;
        RECT 1.1880 1.1410 1.2440 1.5570 ;
    END
    ANTENNADIFFAREA 0.3976 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7940 2.2070 1.1460 2.2630 ;
        RECT 1.0020 2.2630 1.1460 2.3400 ;
        RECT 1.0020 2.2060 1.1460 2.2070 ;
    END
    ANTENNAGATEAREA 0.0165 ;
  END A
  OBS
    LAYER NWELL ;
      RECT -0.1150 3.2240 2.2430 3.4590 ;
      RECT -0.1150 2.3510 0.1150 3.2240 ;
      RECT 2.0130 2.3510 2.2430 3.2240 ;
      RECT 0.5750 2.2340 1.4250 2.7640 ;
      RECT -0.1150 -0.1150 2.2430 0.9930 ;
    LAYER M1 ;
      RECT 0.7750 0.9790 1.4890 1.0350 ;
      RECT 0.7750 1.0350 0.8310 1.0810 ;
      RECT 0.7750 0.9140 0.8310 0.9790 ;
      RECT 0.7390 1.0810 0.8310 1.0820 ;
      RECT 0.7330 0.8580 0.8310 0.9140 ;
      RECT 0.7350 1.0820 0.8310 1.1370 ;
      RECT 0.7330 0.1310 0.7890 0.8580 ;
      RECT 0.7350 1.1370 0.7910 1.5620 ;
      RECT 0.4820 0.9670 0.7250 1.0230 ;
      RECT 0.4820 1.0230 0.5380 1.0910 ;
      RECT 0.4820 0.9090 0.5380 0.9670 ;
      RECT 0.4280 0.8530 0.5380 0.9090 ;
      RECT 0.4300 1.0910 0.5380 1.1380 ;
      RECT 0.4300 1.1380 0.5300 1.1470 ;
      RECT 0.4300 1.1470 0.4860 1.4430 ;
      RECT 0.4280 0.2190 0.4840 0.8530 ;
      RECT 0.1860 0.9670 0.4210 1.0230 ;
      RECT 0.7320 2.3710 0.7880 2.6410 ;
      RECT 0.6400 2.3150 0.7880 2.3710 ;
      RECT 0.6400 2.0790 0.7890 2.1350 ;
      RECT 0.7320 1.8360 0.7880 2.0790 ;
      RECT 0.6400 2.2620 0.6960 2.3150 ;
      RECT 0.3390 2.2060 0.6960 2.2620 ;
      RECT 0.6400 2.1350 0.6960 2.2060 ;
    LAYER PO ;
      RECT 1.7330 0.0690 1.7630 2.7800 ;
      RECT 0.3650 0.0890 0.3950 2.7800 ;
      RECT 1.1250 0.0530 1.1550 2.7780 ;
      RECT 1.8850 0.0690 1.9150 2.7800 ;
      RECT 1.5810 0.0690 1.6110 2.7800 ;
      RECT 1.2770 0.0530 1.3070 2.7800 ;
      RECT 1.4290 0.0530 1.4590 2.7800 ;
      RECT 2.0370 0.0740 2.0670 2.7800 ;
      RECT 0.9730 0.0530 1.0030 2.7800 ;
      RECT 0.8210 0.0780 0.8510 2.7800 ;
      RECT 0.0610 0.0890 0.0910 2.7800 ;
      RECT 0.6690 0.0680 0.6990 2.7810 ;
      RECT 0.5170 0.0890 0.5470 2.7800 ;
      RECT 0.2130 0.0890 0.2430 2.7800 ;
  END
END LSDNX4_LVT

MACRO LSDNX8_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.736 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 3.0100 2.7360 3.0700 ;
        RECT 1.7700 3.0700 1.8800 3.1430 ;
        RECT 1.7700 2.9360 1.8800 3.0100 ;
        RECT 0.8830 2.3430 0.9390 3.0100 ;
        RECT 1.1910 2.5200 1.2410 3.0100 ;
    END
  END VDDH

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.7360 0.0300 ;
        RECT 0.2760 0.0300 0.3320 0.7690 ;
        RECT 2.4040 0.0300 2.4600 0.4670 ;
        RECT 2.1000 0.0300 2.1560 0.7840 ;
        RECT 1.7960 0.0300 1.8520 0.7820 ;
        RECT 1.4920 0.0300 1.5480 0.7750 ;
        RECT 0.5800 0.0300 0.6360 0.8370 ;
        RECT 0.8840 0.0300 0.9400 0.7580 ;
        RECT 1.1880 0.0300 1.2440 0.7750 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 2.7360 3.3740 ;
    END
  END VDDL

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.7360 1.7020 ;
        RECT 0.2500 1.7020 0.3600 1.7750 ;
        RECT 0.2500 1.5680 0.3600 1.6420 ;
        RECT 2.4040 1.2200 2.4600 1.6420 ;
        RECT 1.1880 1.1930 1.2440 1.6420 ;
        RECT 1.4920 1.1930 1.5480 1.6420 ;
        RECT 1.7960 1.1930 1.8520 1.6420 ;
        RECT 2.1000 1.1930 2.1560 1.6420 ;
        RECT 0.8840 1.2500 0.9400 1.6420 ;
        RECT 0.5800 1.1750 0.6360 1.6420 ;
        RECT 0.8840 1.7020 0.9400 2.0250 ;
        RECT 0.2760 1.3050 0.3320 1.5680 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0390 1.0780 2.3450 1.1280 ;
        RECT 1.0390 1.1280 1.0890 1.5620 ;
        RECT 2.2550 1.1280 2.3050 1.5640 ;
        RECT 1.9510 1.1280 2.0010 1.5650 ;
        RECT 1.6470 1.1280 1.6970 1.5650 ;
        RECT 1.3430 1.1280 1.3930 1.5640 ;
        RECT 2.2950 0.9880 2.3450 1.0780 ;
        RECT 2.2950 0.9030 2.4870 0.9880 ;
        RECT 1.0390 0.8540 2.4870 0.9030 ;
        RECT 1.0390 0.8530 2.3450 0.8540 ;
        RECT 1.0390 0.0970 1.0890 0.8530 ;
        RECT 2.2550 0.1090 2.3050 0.8530 ;
        RECT 1.9510 0.0980 2.0010 0.8530 ;
        RECT 1.6470 0.0980 1.6970 0.8530 ;
        RECT 1.3430 0.0980 1.3930 0.8530 ;
    END
    ANTENNADIFFAREA 0.6915 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7940 2.2070 1.1390 2.2630 ;
        RECT 0.9950 2.2630 1.1390 2.3410 ;
    END
    ANTENNAGATEAREA 0.0132 ;
  END A
  OBS
    LAYER NWELL ;
      RECT -0.1150 3.2240 2.8510 3.4590 ;
      RECT 2.4690 2.3510 2.8510 3.2240 ;
      RECT -0.1150 2.3510 0.1150 3.2240 ;
      RECT 0.5750 2.2340 1.4250 2.7640 ;
      RECT -0.1150 -0.1150 2.8510 0.9930 ;
    LAYER M1 ;
      RECT 0.4720 0.9670 0.8770 1.0230 ;
      RECT 0.4720 1.0230 0.5280 1.0910 ;
      RECT 0.4720 0.9090 0.5280 0.9670 ;
      RECT 0.4300 1.0910 0.5280 1.1470 ;
      RECT 0.4280 0.8530 0.5280 0.9090 ;
      RECT 0.4300 1.1470 0.4860 1.4430 ;
      RECT 0.4280 0.2880 0.4840 0.8530 ;
      RECT 0.1860 0.9670 0.4210 1.0230 ;
      RECT 0.9300 0.9670 2.2450 1.0230 ;
      RECT 0.7320 1.1320 0.7880 1.5780 ;
      RECT 0.7320 0.1110 0.7880 0.8480 ;
      RECT 0.9300 1.0230 0.9860 1.0760 ;
      RECT 0.9300 0.9040 0.9860 0.9670 ;
      RECT 0.7320 1.0760 0.9860 1.1320 ;
      RECT 0.7320 0.8480 0.9860 0.9040 ;
      RECT 0.7310 2.3710 0.7870 2.6410 ;
      RECT 0.6390 2.3150 0.7870 2.3710 ;
      RECT 0.6390 2.0790 0.7880 2.1350 ;
      RECT 0.7320 1.9030 0.7880 2.0790 ;
      RECT 0.6390 2.2620 0.6950 2.3150 ;
      RECT 0.3390 2.2060 0.6950 2.2620 ;
      RECT 0.6390 2.1350 0.6950 2.2060 ;
    LAYER PO ;
      RECT 2.6450 0.0740 2.6750 2.7800 ;
      RECT 2.3410 0.0690 2.3710 2.7800 ;
      RECT 1.7330 0.0680 1.7630 2.7800 ;
      RECT 0.3650 0.0890 0.3950 2.7800 ;
      RECT 2.4930 0.0740 2.5230 2.7800 ;
      RECT 1.1250 0.0680 1.1550 2.7780 ;
      RECT 0.8210 0.0680 0.8510 1.6420 ;
      RECT 0.8210 1.7430 0.8510 2.7800 ;
      RECT 1.8850 0.0680 1.9150 2.7800 ;
      RECT 1.5810 0.0680 1.6110 2.7800 ;
      RECT 1.2770 0.0680 1.3070 2.7800 ;
      RECT 1.4290 0.0680 1.4590 2.7800 ;
      RECT 2.0370 0.0680 2.0670 2.7800 ;
      RECT 0.9730 0.0680 1.0030 2.7800 ;
      RECT 2.1890 0.0680 2.2190 2.7800 ;
      RECT 0.0610 0.0890 0.0910 2.7800 ;
      RECT 0.6690 0.0680 0.6990 2.7810 ;
      RECT 0.5170 0.0890 0.5470 2.7800 ;
      RECT 0.2130 0.0890 0.2430 2.7800 ;
  END
END LSDNX8_LVT

MACRO LSUPENCLX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.128 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2460 0.8500 1.4370 0.9840 ;
    END
    ANTENNAGATEAREA 0.0252 ;
  END EN

  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.1280 0.0300 ;
        RECT 1.3430 0.0300 1.3930 0.4130 ;
        RECT 1.7990 0.0300 1.8490 0.4850 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 2.1280 3.3740 ;
    END
  END VDDH

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 3.0100 2.1280 3.0700 ;
        RECT 0.4020 3.0700 0.5120 3.1430 ;
        RECT 0.4020 2.9360 0.5120 3.0100 ;
        RECT 1.1910 2.5200 1.2410 3.0100 ;
        RECT 0.8870 2.5250 0.9370 3.0100 ;
    END
  END VDDL

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.1280 1.7020 ;
        RECT 0.2500 1.7020 0.3600 1.7750 ;
        RECT 0.2500 1.5680 0.3600 1.6420 ;
        RECT 1.4950 1.3070 1.5450 1.6420 ;
        RECT 0.7350 1.7020 0.7850 2.0200 ;
        RECT 0.8870 1.3040 0.9370 1.6420 ;
        RECT 1.7990 1.3030 1.8490 1.6420 ;
        RECT 1.3430 1.7020 1.3930 1.7050 ;
        RECT 1.3430 1.3070 1.3930 1.6420 ;
        RECT 1.0390 1.7020 1.0890 2.0200 ;
        RECT 0.7350 1.3070 0.7850 1.6420 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6870 0.8080 1.7370 0.8420 ;
        RECT 1.6870 0.8420 1.8790 0.9760 ;
        RECT 1.6470 0.7580 1.7370 0.8080 ;
        RECT 1.6870 0.9760 1.7370 1.1770 ;
        RECT 1.6470 0.2110 1.6970 0.7580 ;
        RECT 1.1910 1.1770 1.7370 1.2270 ;
        RECT 1.6470 1.2270 1.6970 1.5870 ;
        RECT 1.1910 1.2270 1.2410 1.5870 ;
    END
    ANTENNADIFFAREA 0.1672 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7940 2.2130 1.1600 2.2630 ;
        RECT 0.9970 2.2630 1.1600 2.3650 ;
    END
    ANTENNAGATEAREA 0.0468 ;
  END A
  OBS
    LAYER NWELL ;
      RECT -0.1150 3.2240 2.2430 3.4590 ;
      RECT -0.1150 2.3510 0.1150 3.2240 ;
      RECT 2.0130 2.3510 2.2430 3.2240 ;
      RECT 0.5750 2.2340 1.4250 2.7640 ;
      RECT -0.1150 -0.1150 2.2430 0.9930 ;
    LAYER M1 ;
      RECT 1.1910 0.5270 1.5450 0.5770 ;
      RECT 1.4950 0.1520 1.5450 0.5270 ;
      RECT 1.1910 0.1640 1.2410 0.5270 ;
      RECT 0.8870 0.1140 1.2410 0.1640 ;
      RECT 0.8870 0.1640 0.9370 0.1790 ;
      RECT 0.7360 0.1790 0.9370 0.2040 ;
      RECT 0.7350 0.2040 0.9370 0.2290 ;
      RECT 0.7350 0.2290 0.7850 0.4130 ;
      RECT 0.8870 0.2290 0.9370 0.4240 ;
      RECT 1.5710 1.0100 1.6210 1.0380 ;
      RECT 1.0390 1.0380 1.6210 1.0880 ;
      RECT 1.5710 1.0880 1.6210 1.1160 ;
      RECT 1.0390 1.0880 1.0890 1.5870 ;
      RECT 1.0390 1.0140 1.1290 1.0380 ;
      RECT 1.0790 0.9110 1.1290 1.0140 ;
      RECT 0.6430 0.8610 1.1290 0.9110 ;
      RECT 1.0790 0.5770 1.1290 0.8610 ;
      RECT 1.0390 0.5160 1.1290 0.5770 ;
      RECT 1.0390 0.2740 1.0890 0.5160 ;
      RECT 0.5430 0.6910 1.0290 0.7410 ;
      RECT 0.5430 0.6840 0.6330 0.6910 ;
      RECT 0.5430 0.7410 0.5930 1.2960 ;
      RECT 0.5830 0.2300 0.6330 0.6840 ;
      RECT 0.5430 1.2960 0.6330 1.3460 ;
      RECT 0.5830 1.3460 0.6330 1.5870 ;
      RECT 1.0390 2.4730 1.0890 2.6900 ;
      RECT 0.6590 2.4230 1.0890 2.4730 ;
      RECT 0.6590 2.1330 0.7090 2.4230 ;
      RECT 0.6590 2.0830 0.9370 2.1330 ;
      RECT 0.8870 1.8670 0.9370 2.0830 ;
      RECT 0.7350 2.4730 0.7850 2.6900 ;
    LAYER PO ;
      RECT 1.7330 0.0690 1.7630 2.7800 ;
      RECT 0.3650 0.0890 0.3950 2.7800 ;
      RECT 1.5810 0.0640 1.6110 1.6690 ;
      RECT 1.1250 0.0870 1.1550 2.7780 ;
      RECT 0.9730 0.0890 1.0030 1.0250 ;
      RECT 1.8850 0.0690 1.9150 2.7800 ;
      RECT 0.8210 1.7710 0.8510 2.7820 ;
      RECT 0.9730 1.1630 1.0030 2.7820 ;
      RECT 1.2770 0.0750 1.3070 2.7800 ;
      RECT 1.4290 0.0750 1.4590 2.7800 ;
      RECT 2.0370 0.0740 2.0670 2.7800 ;
      RECT 0.6690 0.0890 0.6990 1.0250 ;
      RECT 0.8210 0.0780 0.8510 1.6700 ;
      RECT 0.0610 0.0890 0.0910 2.7800 ;
      RECT 0.6690 1.1780 0.6990 2.7810 ;
      RECT 0.5170 0.0890 0.5470 2.7800 ;
      RECT 0.2130 0.0890 0.2430 2.7800 ;
  END
END LSUPENCLX1_LVT

MACRO LSUPENCLX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.128 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9420 0.8500 1.1330 0.9840 ;
    END
    ANTENNAGATEAREA 0.0324 ;
  END EN

  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.1280 0.0300 ;
        RECT 1.0390 0.0300 1.0890 0.4130 ;
        RECT 1.7990 0.0300 1.8490 0.4850 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 2.1280 3.3740 ;
    END
  END VDDH

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 3.0100 2.1280 3.0700 ;
        RECT 1.7700 3.0700 1.8800 3.1430 ;
        RECT 1.7700 2.9360 1.8800 3.0100 ;
        RECT 1.1910 2.5200 1.2410 3.0100 ;
        RECT 0.9110 2.7350 0.9610 3.0100 ;
        RECT 0.8870 2.6740 0.9610 2.7350 ;
        RECT 0.8870 2.5250 0.9370 2.6740 ;
    END
  END VDDL

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.1280 1.7020 ;
        RECT 1.7700 1.7020 1.8800 1.7750 ;
        RECT 1.7700 1.5680 1.8800 1.6420 ;
        RECT 1.4950 1.4110 1.5450 1.6420 ;
        RECT 0.7350 1.7020 0.7850 2.0200 ;
        RECT 0.5830 1.3540 0.6330 1.6420 ;
        RECT 1.0390 1.3620 1.0890 1.6420 ;
        RECT 1.0390 1.7020 1.0890 2.0200 ;
        RECT 0.4310 1.3620 0.4810 1.6420 ;
        RECT 1.7990 1.3030 1.8490 1.5680 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6470 0.2110 1.6970 0.4960 ;
        RECT 1.6470 0.4960 1.7370 0.5460 ;
        RECT 1.6870 0.5460 1.7370 0.8160 ;
        RECT 1.3430 0.8160 1.7370 0.8420 ;
        RECT 1.3430 0.6470 1.3930 0.8160 ;
        RECT 1.3430 0.8420 1.8790 0.8660 ;
        RECT 1.6870 0.8660 1.8790 0.9760 ;
        RECT 1.6870 0.9760 1.7370 1.1770 ;
        RECT 0.8870 1.1770 1.7370 1.2270 ;
        RECT 1.1910 1.2270 1.2410 1.5870 ;
        RECT 1.3430 1.2270 1.3930 1.5870 ;
        RECT 0.8870 1.2270 0.9370 1.5870 ;
        RECT 1.6870 1.2270 1.7370 1.2990 ;
        RECT 1.6470 1.2990 1.7370 1.3720 ;
        RECT 1.6470 1.3720 1.6970 1.5870 ;
    END
    ANTENNADIFFAREA 0.3038 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7940 2.2130 1.1600 2.2630 ;
        RECT 0.9970 2.2630 1.1600 2.3650 ;
    END
    ANTENNAGATEAREA 0.0489 ;
  END A
  OBS
    LAYER NWELL ;
      RECT -0.1150 3.2240 2.2430 3.4590 ;
      RECT -0.1150 2.3510 0.1150 3.2240 ;
      RECT 2.0130 2.3510 2.2430 3.2240 ;
      RECT 0.5750 2.2340 1.4250 2.7640 ;
      RECT -0.1150 -0.1150 2.2430 0.9930 ;
    LAYER M1 ;
      RECT 1.1150 0.6950 1.1650 0.7170 ;
      RECT 0.9460 0.7170 1.1650 0.7670 ;
      RECT 1.1150 0.7670 1.1650 0.7830 ;
      RECT 0.8110 2.8400 0.8610 2.8620 ;
      RECT 0.6420 2.8620 0.8610 2.9120 ;
      RECT 0.8110 2.9120 0.8610 2.9280 ;
      RECT 0.8870 0.4960 1.5450 0.5460 ;
      RECT 1.1910 0.1880 1.2410 0.4960 ;
      RECT 1.4950 0.1520 1.5450 0.4960 ;
      RECT 0.8870 0.1640 0.9370 0.4960 ;
      RECT 0.5830 0.1140 0.9400 0.1640 ;
      RECT 0.5830 0.1640 0.6330 0.1790 ;
      RECT 0.4320 0.1790 0.6330 0.2040 ;
      RECT 0.4310 0.2040 0.6330 0.2290 ;
      RECT 0.4310 0.2290 0.4810 0.4130 ;
      RECT 0.5830 0.2290 0.6330 0.4240 ;
      RECT 1.5710 1.0100 1.6210 1.0380 ;
      RECT 0.7350 1.0380 1.6210 1.0880 ;
      RECT 1.5710 1.0880 1.6210 1.1160 ;
      RECT 0.7350 1.0880 0.7850 1.5870 ;
      RECT 0.7350 1.0140 0.8250 1.0380 ;
      RECT 0.7750 0.8600 0.8250 1.0140 ;
      RECT 0.3390 0.8100 0.8250 0.8600 ;
      RECT 0.7750 0.5770 0.8250 0.8100 ;
      RECT 0.7350 0.5160 0.8250 0.5770 ;
      RECT 0.7350 0.2740 0.7850 0.5160 ;
      RECT 0.2390 0.6910 0.7250 0.7410 ;
      RECT 0.2390 0.6840 0.3290 0.6910 ;
      RECT 0.2390 0.7410 0.2890 1.2990 ;
      RECT 0.2790 0.2300 0.3290 0.6840 ;
      RECT 0.2390 1.2990 0.3290 1.3650 ;
      RECT 0.2790 1.3650 0.3290 1.5870 ;
      RECT 0.6590 2.4230 1.0890 2.4730 ;
      RECT 1.0390 2.4730 1.0890 2.6900 ;
      RECT 0.6590 2.2630 0.7090 2.4230 ;
      RECT 0.3310 2.2130 0.7090 2.2630 ;
      RECT 0.6590 2.1330 0.7090 2.2130 ;
      RECT 0.6590 2.0830 0.9370 2.1330 ;
      RECT 0.8870 1.8670 0.9370 2.0830 ;
      RECT 0.7350 2.4730 0.7850 2.6900 ;
    LAYER PO ;
      RECT 1.7330 0.0690 1.7630 2.7800 ;
      RECT 0.3650 1.1290 0.3950 2.7800 ;
      RECT 1.5810 0.0650 1.6110 1.6690 ;
      RECT 0.8210 0.0860 0.8510 1.6470 ;
      RECT 1.1250 0.0870 1.1550 2.7780 ;
      RECT 0.6690 0.0890 0.6990 0.9140 ;
      RECT 1.8850 0.0690 1.9150 2.7800 ;
      RECT 0.8210 1.8120 0.8510 2.9270 ;
      RECT 0.9730 0.0860 1.0030 1.6680 ;
      RECT 1.2770 0.0750 1.3070 2.7800 ;
      RECT 1.4290 0.0640 1.4590 2.7170 ;
      RECT 2.0370 0.0740 2.0670 2.7800 ;
      RECT 0.3650 0.0870 0.3950 0.9090 ;
      RECT 0.9730 1.7690 1.0030 2.7820 ;
      RECT 0.6690 1.1350 0.6990 2.9230 ;
      RECT 0.5170 0.0780 0.5470 2.7800 ;
      RECT 0.2130 0.0890 0.2430 2.7800 ;
      RECT 0.0610 0.0890 0.0910 2.7800 ;
  END
END LSUPENCLX2_LVT

MACRO LSUPENCLX4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.04 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9420 0.8500 1.1330 0.9840 ;
    END
    ANTENNAGATEAREA 0.0402 ;
  END EN

  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.0400 0.0300 ;
        RECT 1.0390 0.0300 1.0890 0.4130 ;
        RECT 2.7110 0.0300 2.7610 0.4850 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 3.0400 3.3740 ;
    END
  END VDDH

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 3.0100 3.0400 3.0700 ;
        RECT 1.7700 3.0700 1.8800 3.1430 ;
        RECT 1.7700 2.9360 1.8800 3.0100 ;
        RECT 1.1910 2.5200 1.2410 3.0100 ;
        RECT 0.9110 2.7350 0.9610 3.0100 ;
        RECT 0.8870 2.6740 0.9610 2.7350 ;
        RECT 0.8870 2.5250 0.9370 2.6740 ;
    END
  END VDDL

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.0400 1.7020 ;
        RECT 2.6820 1.7020 2.7920 1.7750 ;
        RECT 2.6820 1.5680 2.7920 1.6420 ;
        RECT 0.5830 1.3200 0.6330 1.6420 ;
        RECT 1.0390 1.7020 1.0890 1.7050 ;
        RECT 1.0390 1.3620 1.0890 1.6420 ;
        RECT 0.4310 1.3280 0.4810 1.6420 ;
        RECT 2.4070 1.4110 2.4570 1.6420 ;
        RECT 2.1030 1.4110 2.1530 1.6420 ;
        RECT 1.6470 1.2970 1.6970 1.6420 ;
        RECT 0.7350 1.7020 0.7850 2.0200 ;
        RECT 1.3430 1.4090 1.3930 1.6420 ;
        RECT 2.7110 1.3030 2.7610 1.5680 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5830 0.9940 2.8190 1.1280 ;
        RECT 2.5830 0.8690 2.6330 0.9940 ;
        RECT 2.5830 1.1280 2.6330 1.2880 ;
        RECT 1.9510 0.8200 2.6330 0.8690 ;
        RECT 1.9510 1.2880 2.6330 1.3380 ;
        RECT 1.9510 0.8190 2.6320 0.8200 ;
        RECT 2.2550 1.3380 2.3050 1.5840 ;
        RECT 1.9510 1.3380 2.0010 1.5840 ;
        RECT 2.5590 1.3380 2.6330 1.3680 ;
        RECT 2.5590 0.3040 2.6090 0.8190 ;
        RECT 2.2550 0.2140 2.3050 0.8190 ;
        RECT 1.9510 0.3040 2.0010 0.8190 ;
        RECT 2.5590 1.3680 2.6090 1.5840 ;
    END
    ANTENNADIFFAREA 0.4526 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7940 2.2130 1.1600 2.2630 ;
        RECT 0.9970 2.2630 1.1600 2.3650 ;
    END
    ANTENNAGATEAREA 0.0234 ;
  END A
  OBS
    LAYER NWELL ;
      RECT -0.1150 3.2240 3.1550 3.4590 ;
      RECT -0.1150 2.3510 0.1150 3.2240 ;
      RECT 2.9250 2.3510 3.1550 3.2240 ;
      RECT 0.5750 2.2340 1.4250 2.7640 ;
      RECT -0.1150 -0.1150 3.1550 0.9930 ;
    LAYER M1 ;
      RECT 1.8390 1.0380 2.5330 1.0880 ;
      RECT 2.4830 1.0880 2.5330 1.1230 ;
      RECT 2.4830 0.9980 2.5330 1.0380 ;
      RECT 1.8390 0.8080 1.8890 1.0380 ;
      RECT 1.8390 1.0880 1.8890 1.2720 ;
      RECT 1.7990 0.7820 1.8890 0.8080 ;
      RECT 1.7990 1.2720 1.8890 1.3220 ;
      RECT 1.7990 0.7580 1.8880 0.7820 ;
      RECT 1.7990 1.3220 1.8490 1.5840 ;
      RECT 1.7990 0.2140 1.8490 0.7580 ;
      RECT 2.4070 0.1400 2.4570 0.7630 ;
      RECT 1.3430 0.0900 2.4570 0.1400 ;
      RECT 1.6470 0.1400 1.6970 0.7970 ;
      RECT 1.3430 0.1400 1.3930 0.4960 ;
      RECT 0.8870 0.4960 1.3930 0.5460 ;
      RECT 1.1910 0.1880 1.2410 0.4960 ;
      RECT 0.8870 0.1640 0.9370 0.4960 ;
      RECT 0.5830 0.1140 0.9400 0.1640 ;
      RECT 0.5830 0.1640 0.6330 0.1790 ;
      RECT 0.4320 0.1790 0.6330 0.1970 ;
      RECT 0.4310 0.1970 0.6330 0.2290 ;
      RECT 0.5830 0.2290 0.6330 0.4410 ;
      RECT 0.4310 0.2290 0.4810 0.4310 ;
      RECT 2.1030 0.1400 2.1530 0.7630 ;
      RECT 1.1150 0.6950 1.1650 0.7170 ;
      RECT 0.9460 0.7170 1.1650 0.7670 ;
      RECT 1.1150 0.7670 1.1650 0.7830 ;
      RECT 0.8110 2.8400 0.8610 2.8620 ;
      RECT 0.6420 2.8620 0.8610 2.9120 ;
      RECT 0.8110 2.9120 0.8610 2.9280 ;
      RECT 1.7230 1.0680 1.7730 1.1420 ;
      RECT 1.5350 1.0180 1.7730 1.0680 ;
      RECT 1.5350 1.0680 1.5850 1.1770 ;
      RECT 1.5350 0.5650 1.5850 1.0180 ;
      RECT 1.4950 1.1770 1.5850 1.2500 ;
      RECT 1.4950 0.5150 1.5850 0.5650 ;
      RECT 1.4950 1.2500 1.5450 1.5840 ;
      RECT 1.4950 0.2280 1.5450 0.5150 ;
      RECT 0.7350 1.0380 1.4690 1.0880 ;
      RECT 1.4190 0.7830 1.4690 1.0380 ;
      RECT 0.7350 1.0880 0.7850 1.5840 ;
      RECT 0.7350 1.0140 0.8250 1.0380 ;
      RECT 0.7750 0.9110 0.8250 1.0140 ;
      RECT 0.3390 0.8610 0.8250 0.9110 ;
      RECT 0.7750 0.5770 0.8250 0.8610 ;
      RECT 0.7350 0.5160 0.8250 0.5770 ;
      RECT 0.7350 0.2740 0.7850 0.5160 ;
      RECT 0.2390 0.6910 0.7250 0.7410 ;
      RECT 0.2390 0.6840 0.3290 0.6910 ;
      RECT 0.2390 0.7410 0.2890 1.2960 ;
      RECT 0.2790 0.2300 0.3290 0.6840 ;
      RECT 0.2390 1.2960 0.3290 1.3460 ;
      RECT 0.2790 1.3460 0.3290 1.5840 ;
      RECT 0.8870 1.8670 0.9370 2.0830 ;
      RECT 0.6590 2.0830 0.9370 2.1330 ;
      RECT 0.6590 2.4230 0.7850 2.4730 ;
      RECT 0.7350 2.4730 0.7850 2.6900 ;
      RECT 0.6590 2.1330 0.7090 2.2130 ;
      RECT 0.3310 2.2130 0.7090 2.2630 ;
      RECT 0.6590 2.2630 0.7090 2.4230 ;
      RECT 0.8870 1.1770 1.3460 1.2270 ;
      RECT 0.8870 1.2270 0.9370 1.5840 ;
      RECT 1.1910 1.2270 1.2410 1.5840 ;
      RECT 1.2350 1.9510 2.7050 2.0010 ;
    LAYER PO ;
      RECT 0.3650 0.0870 0.3950 0.9280 ;
      RECT 0.9730 1.7690 1.0030 2.7820 ;
      RECT 0.6690 1.1350 0.6990 2.9230 ;
      RECT 0.5170 0.0780 0.5470 2.7800 ;
      RECT 0.2130 0.0890 0.2430 2.7800 ;
      RECT 0.0610 0.0890 0.0910 2.7800 ;
      RECT 2.7970 0.0680 2.8270 2.7800 ;
      RECT 2.9490 0.0670 2.9790 2.7800 ;
      RECT 1.7330 0.0670 1.7630 2.7800 ;
      RECT 2.3410 0.0680 2.3710 2.7800 ;
      RECT 2.1890 0.0680 2.2190 2.7800 ;
      RECT 2.4930 0.0670 2.5230 2.7800 ;
      RECT 2.6450 0.0680 2.6750 2.7800 ;
      RECT 0.3650 1.1290 0.3950 2.7800 ;
      RECT 1.5810 0.0690 1.6110 2.7800 ;
      RECT 0.8210 0.0860 0.8510 1.6470 ;
      RECT 1.1250 0.0870 1.1550 2.7780 ;
      RECT 0.6690 0.0890 0.6990 0.8640 ;
      RECT 1.8850 0.0680 1.9150 2.7800 ;
      RECT 0.8210 1.8120 0.8510 2.9270 ;
      RECT 1.4290 0.0750 1.4590 2.7800 ;
      RECT 0.9730 0.0860 1.0030 1.6680 ;
      RECT 1.2770 0.0750 1.3070 2.7800 ;
      RECT 2.0370 0.0680 2.0670 2.7800 ;
  END
END LSUPENCLX4_LVT

MACRO LSUPENCLX8_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.712 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.2550 1.0090 4.4660 1.1300 ;
        RECT 4.2550 0.8680 4.3050 1.0090 ;
        RECT 4.2550 1.1300 4.3050 1.2880 ;
        RECT 3.0150 0.8180 4.3050 0.8680 ;
        RECT 3.0150 1.2880 4.3050 1.3380 ;
        RECT 3.9270 0.2130 3.9770 0.8180 ;
        RECT 3.6230 0.2130 3.6730 0.8180 ;
        RECT 3.3190 0.2130 3.3690 0.8180 ;
        RECT 3.0150 0.2110 3.0650 0.8180 ;
        RECT 4.2310 0.7730 4.3050 0.8180 ;
        RECT 3.9270 1.3380 3.9770 1.5840 ;
        RECT 3.6230 1.3380 3.6730 1.5840 ;
        RECT 3.3190 1.3380 3.3690 1.5840 ;
        RECT 3.0150 1.3380 3.0650 1.5840 ;
        RECT 4.2310 1.3380 4.3050 1.4140 ;
        RECT 4.2310 0.2110 4.2810 0.7730 ;
        RECT 4.2310 1.4140 4.2810 1.5840 ;
    END
    ANTENNADIFFAREA 0.9344 ;
  END Y

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0060 1.9080 2.1970 2.0420 ;
    END
    ANTENNAGATEAREA 0.2928 ;
  END EN

  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.7120 0.0300 ;
        RECT 1.9510 0.0300 2.0010 0.7430 ;
        RECT 1.6470 0.0300 1.6970 0.7430 ;
        RECT 1.3430 0.0300 1.3930 0.7430 ;
        RECT 1.0390 0.0300 1.0890 0.7430 ;
        RECT 4.3830 0.0300 4.4330 0.4360 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 4.7120 3.3740 ;
    END
  END VDDH

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 3.0100 4.7120 3.0700 ;
        RECT 2.9860 3.0700 3.0960 3.1430 ;
        RECT 2.9860 2.9360 3.0960 3.0100 ;
        RECT 1.1910 2.5200 1.2410 3.0100 ;
        RECT 0.9110 2.7350 0.9610 3.0100 ;
        RECT 0.8870 2.6740 0.9610 2.7350 ;
        RECT 0.8870 2.5250 0.9370 2.6740 ;
    END
  END VDDL

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.7120 1.7020 ;
        RECT 0.4020 1.7020 0.5120 1.7750 ;
        RECT 0.4020 1.5680 0.5120 1.6420 ;
        RECT 3.4710 1.4110 3.5210 1.6420 ;
        RECT 3.1670 1.4110 3.2170 1.6420 ;
        RECT 2.7110 1.4110 2.7610 1.6420 ;
        RECT 0.7350 1.7020 0.7850 2.0200 ;
        RECT 2.2550 1.3980 2.3050 1.6420 ;
        RECT 0.5830 1.2360 0.6330 1.6420 ;
        RECT 4.3830 1.3030 4.4330 1.6420 ;
        RECT 1.0390 1.4040 1.0890 1.6420 ;
        RECT 1.0390 1.7020 1.0890 2.0200 ;
        RECT 1.6470 1.7020 1.6970 1.7050 ;
        RECT 1.6470 1.4000 1.6970 1.6420 ;
        RECT 1.3430 1.7020 1.3930 1.7050 ;
        RECT 1.3430 1.4050 1.3930 1.6420 ;
        RECT 1.9510 1.7020 2.0010 1.7050 ;
        RECT 1.9510 1.4020 2.0010 1.6420 ;
        RECT 4.0790 1.4110 4.1290 1.6420 ;
        RECT 3.7750 1.4110 3.8250 1.6420 ;
        RECT 0.4310 1.2360 0.4810 1.5680 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7940 2.2130 1.1600 2.2630 ;
        RECT 0.9970 2.2630 1.1600 2.3650 ;
    END
    ANTENNAGATEAREA 0.0486 ;
  END A
  OBS
    LAYER NWELL ;
      RECT -0.1150 3.2240 4.8270 3.4590 ;
      RECT -0.1150 2.3510 0.1150 3.2240 ;
      RECT 4.5970 2.3510 4.8270 3.2240 ;
      RECT 0.5750 2.2340 1.4250 2.7640 ;
      RECT -0.1150 -0.1150 4.8270 0.9930 ;
    LAYER M1 ;
      RECT 0.2390 0.6910 0.7250 0.7410 ;
      RECT 0.2790 1.3300 0.3290 1.5840 ;
      RECT 0.2390 1.2800 0.3290 1.3300 ;
      RECT 0.2390 0.7410 0.2890 1.2800 ;
      RECT 0.2390 0.6840 0.3290 0.6910 ;
      RECT 0.2790 0.2300 0.3290 0.6840 ;
      RECT 0.6590 2.4230 1.0890 2.4730 ;
      RECT 1.0390 2.4730 1.0890 2.6900 ;
      RECT 0.6590 2.2630 0.7090 2.4230 ;
      RECT 0.3310 2.2130 0.7090 2.2630 ;
      RECT 0.6590 2.1330 0.7090 2.2130 ;
      RECT 0.6590 2.0830 0.9370 2.1330 ;
      RECT 0.8870 1.8670 0.9370 2.0830 ;
      RECT 0.7350 2.4730 0.7850 2.6900 ;
      RECT 2.1460 1.7890 4.4080 1.8390 ;
      RECT 2.1790 1.0740 2.2290 1.2500 ;
      RECT 0.8870 1.2500 2.2290 1.3000 ;
      RECT 0.8870 1.3000 0.9370 1.5840 ;
      RECT 1.1910 1.3000 1.2410 1.5840 ;
      RECT 1.4950 1.3000 1.5450 1.5840 ;
      RECT 1.7990 1.3000 1.8490 1.5840 ;
      RECT 2.1030 1.3000 2.1530 1.5840 ;
      RECT 4.0790 0.1390 4.1290 0.7620 ;
      RECT 2.2550 0.1380 4.1290 0.1390 ;
      RECT 2.1030 0.0890 4.1290 0.1380 ;
      RECT 2.2550 0.1390 2.3050 0.7310 ;
      RECT 2.7110 0.1390 2.7610 0.7590 ;
      RECT 2.1030 0.1380 2.1530 0.8080 ;
      RECT 2.1030 0.0880 2.2830 0.0890 ;
      RECT 0.8870 0.8080 2.1530 0.8580 ;
      RECT 3.1670 0.1390 3.2170 0.7590 ;
      RECT 3.4710 0.1390 3.5210 0.7610 ;
      RECT 3.7750 0.1390 3.8250 0.7310 ;
      RECT 0.8870 0.1380 0.9370 0.8080 ;
      RECT 0.5830 0.0880 0.9370 0.1380 ;
      RECT 0.5830 0.1380 0.6330 0.1790 ;
      RECT 0.4320 0.1790 0.6330 0.2040 ;
      RECT 0.4310 0.2040 0.6330 0.2290 ;
      RECT 0.4310 0.2290 0.4810 0.4130 ;
      RECT 0.5830 0.2290 0.6330 0.4240 ;
      RECT 1.1910 0.1270 1.2410 0.8080 ;
      RECT 1.4950 0.1270 1.5450 0.8080 ;
      RECT 1.7990 0.1270 1.8490 0.8080 ;
      RECT 2.9030 1.0380 4.2050 1.0880 ;
      RECT 4.1550 1.0880 4.2050 1.1230 ;
      RECT 4.1550 0.9220 4.2050 1.0380 ;
      RECT 2.5590 1.3380 2.6090 1.5840 ;
      RECT 2.5590 0.2110 2.6090 0.8180 ;
      RECT 2.9030 1.0880 2.9530 1.2880 ;
      RECT 2.9030 0.8680 2.9530 1.0380 ;
      RECT 2.5590 1.2880 2.9530 1.3380 ;
      RECT 2.5590 0.8180 2.9530 0.8680 ;
      RECT 2.8630 1.3380 2.9530 1.3720 ;
      RECT 2.8630 0.8020 2.9530 0.8180 ;
      RECT 2.8630 1.3720 2.9130 1.5840 ;
      RECT 2.8630 0.2130 2.9130 0.8020 ;
      RECT 0.9360 1.0920 2.0770 1.1420 ;
      RECT 2.0270 1.1420 2.0770 1.1680 ;
      RECT 2.0270 1.0760 2.0770 1.0920 ;
      RECT 0.8110 2.8400 0.8610 2.8620 ;
      RECT 0.6420 2.8620 0.8610 2.9120 ;
      RECT 0.8110 2.9120 0.8610 2.9280 ;
      RECT 2.4470 1.0380 2.8530 1.0880 ;
      RECT 2.4470 0.7650 2.4970 1.0380 ;
      RECT 2.4470 1.0880 2.4970 1.2020 ;
      RECT 2.4070 0.7050 2.4970 0.7650 ;
      RECT 2.4070 1.2020 2.4970 1.2500 ;
      RECT 2.4070 0.2610 2.4570 0.7050 ;
      RECT 2.4070 1.2500 2.4960 1.2520 ;
      RECT 2.4070 1.2520 2.4570 1.5840 ;
      RECT 0.7350 0.9700 2.3810 1.0200 ;
      RECT 2.3310 0.8190 2.3810 0.9700 ;
      RECT 0.7350 1.0200 0.7850 1.5840 ;
      RECT 0.7750 0.8410 0.8250 0.9700 ;
      RECT 0.3390 0.7910 0.8250 0.8410 ;
      RECT 0.7750 0.5770 0.8250 0.7910 ;
      RECT 0.7350 0.5160 0.8250 0.5770 ;
      RECT 0.7350 0.2740 0.7850 0.5160 ;
    LAYER PO ;
      RECT 4.6210 0.0740 4.6510 2.7800 ;
      RECT 4.3170 0.0690 4.3470 2.7800 ;
      RECT 4.4690 0.0740 4.4990 2.7800 ;
      RECT 4.1650 0.0670 4.1950 2.7800 ;
      RECT 4.0130 0.0670 4.0430 2.7800 ;
      RECT 3.7090 0.0670 3.7390 2.7800 ;
      RECT 3.8610 0.0670 3.8910 2.7800 ;
      RECT 3.4050 0.0670 3.4350 2.7800 ;
      RECT 3.5570 0.0670 3.5870 2.7800 ;
      RECT 3.2530 0.0670 3.2830 2.7800 ;
      RECT 3.1010 0.0670 3.1310 2.7800 ;
      RECT 2.7970 0.0670 2.8270 2.7800 ;
      RECT 2.9490 0.0670 2.9790 2.7800 ;
      RECT 2.1890 0.0670 2.2190 2.7800 ;
      RECT 2.3410 0.0670 2.3710 2.7800 ;
      RECT 2.6450 0.0670 2.6750 2.7800 ;
      RECT 1.7330 0.0670 1.7630 2.7800 ;
      RECT 0.3650 1.1280 0.3950 2.7800 ;
      RECT 2.4930 0.0670 2.5230 2.7780 ;
      RECT 0.8210 0.0860 0.8510 1.6470 ;
      RECT 1.1250 0.0670 1.1550 2.7780 ;
      RECT 0.6690 0.0890 0.6990 0.9130 ;
      RECT 1.8850 0.0670 1.9150 2.7800 ;
      RECT 0.8210 1.8120 0.8510 2.9270 ;
      RECT 0.9730 0.0670 1.0030 1.6680 ;
      RECT 1.5810 0.0670 1.6110 2.7800 ;
      RECT 1.2770 0.0670 1.3070 2.7800 ;
      RECT 1.4290 0.0670 1.4590 2.7800 ;
      RECT 2.0370 0.0670 2.0670 2.7800 ;
      RECT 0.3650 0.0870 0.3950 0.9110 ;
      RECT 0.9730 1.7690 1.0030 2.7820 ;
      RECT 0.6690 1.1350 0.6990 2.9230 ;
      RECT 0.5170 0.0780 0.5470 2.7800 ;
      RECT 0.2130 0.0890 0.2430 2.7800 ;
      RECT 0.0610 0.0890 0.0910 2.7800 ;
  END
END LSUPENCLX8_LVT

MACRO LSUPENX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.28 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7690 0.8570 1.8790 0.8870 ;
        RECT 1.6470 0.8870 1.8790 0.9370 ;
        RECT 1.7690 0.9370 1.8790 0.9670 ;
        RECT 1.6470 0.5890 1.6970 0.8870 ;
        RECT 1.7990 0.9670 1.8490 1.5660 ;
        RECT 1.0390 0.5390 1.6970 0.5890 ;
        RECT 1.0390 0.1790 1.0890 0.5390 ;
        RECT 1.0390 0.5890 1.0890 0.9050 ;
        RECT 1.6470 0.1190 1.6970 0.5390 ;
    END
    ANTENNADIFFAREA 0.206 ;
  END Y

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3130 2.2240 1.4950 2.3340 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END EN

  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.2800 0.0300 ;
        RECT 1.4950 0.0300 1.5450 0.4840 ;
        RECT 0.5830 0.0300 0.6330 0.4590 ;
        RECT 0.4310 0.0300 0.4810 0.4640 ;
        RECT 1.7990 0.0300 1.8490 0.7530 ;
        RECT 0.8870 0.0300 0.9370 0.8730 ;
        RECT 1.9510 0.0300 2.0010 0.5260 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 2.2800 3.3740 ;
    END
  END VDDH

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 3.0100 2.2800 3.0700 ;
        RECT 1.6180 3.0700 1.7280 3.1430 ;
        RECT 1.6180 2.9360 1.7280 3.0100 ;
        RECT 1.1910 2.5200 1.2410 3.0100 ;
        RECT 0.9110 2.7350 0.9610 3.0100 ;
        RECT 0.8870 2.6740 0.9610 2.7350 ;
        RECT 0.8870 2.5250 0.9370 2.6740 ;
    END
  END VDDL

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.2800 1.7020 ;
        RECT 1.9220 1.7020 2.0320 1.7750 ;
        RECT 1.9220 1.5680 2.0320 1.6420 ;
        RECT 1.0390 1.3520 1.0890 1.6420 ;
        RECT 1.4950 1.4820 1.5450 1.6420 ;
        RECT 1.9510 1.3030 2.0010 1.5680 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7940 2.2130 1.1600 2.2630 ;
        RECT 0.9970 2.2630 1.1600 2.3650 ;
    END
    ANTENNAGATEAREA 0.0492 ;
  END A
  OBS
    LAYER NWELL ;
      RECT -0.1150 3.2240 2.3950 3.4590 ;
      RECT -0.1150 2.3510 0.1150 3.2240 ;
      RECT 2.1650 2.3510 2.3950 3.2240 ;
      RECT 0.5750 2.2340 1.4250 2.7640 ;
      RECT -0.1150 -0.1150 2.3950 0.9930 ;
    LAYER M1 ;
      RECT 0.2390 0.6920 0.7250 0.7420 ;
      RECT 0.2390 0.7420 0.2890 1.0470 ;
      RECT 0.2390 0.6840 0.3290 0.6920 ;
      RECT 0.2390 1.0470 0.3290 1.0970 ;
      RECT 0.2790 0.2800 0.3290 0.6840 ;
      RECT 0.2790 1.0970 0.3290 1.5820 ;
      RECT 0.8110 2.8400 0.8610 2.8620 ;
      RECT 0.6420 2.8620 0.8610 2.9120 ;
      RECT 0.8110 2.9120 0.8610 2.9280 ;
      RECT 0.9360 1.1020 1.4330 1.1520 ;
      RECT 1.3430 1.1520 1.3930 1.5900 ;
      RECT 1.3830 0.9050 1.4330 1.1020 ;
      RECT 1.3430 0.8550 1.4330 0.9050 ;
      RECT 1.3430 0.6390 1.3930 0.8550 ;
      RECT 0.7350 1.0240 1.3330 1.0510 ;
      RECT 0.7750 1.0010 1.3330 1.0240 ;
      RECT 0.7350 1.0510 0.8250 1.0970 ;
      RECT 0.7750 0.8690 0.8250 1.0010 ;
      RECT 0.7350 1.0970 0.7850 1.4110 ;
      RECT 0.3390 0.8190 0.8250 0.8690 ;
      RECT 0.7750 0.5510 0.8250 0.8190 ;
      RECT 0.7350 0.5010 0.8250 0.5510 ;
      RECT 0.7350 0.2740 0.7850 0.5010 ;
      RECT 1.1910 1.3000 1.2410 1.5870 ;
      RECT 0.8870 1.2500 1.2410 1.3000 ;
      RECT 0.8870 1.3000 0.9370 1.5310 ;
      RECT 0.8870 1.2430 0.9370 1.2500 ;
      RECT 0.4310 1.5310 0.9370 1.5810 ;
      RECT 0.5830 1.2220 0.6330 1.5310 ;
      RECT 0.4310 1.5810 0.4810 1.5820 ;
      RECT 0.4310 1.1540 0.4810 1.5310 ;
      RECT 0.4310 1.1040 0.5730 1.1540 ;
      RECT 1.0390 2.4730 1.0890 2.6900 ;
      RECT 0.6590 2.4230 1.0890 2.4730 ;
      RECT 0.6590 2.2630 0.7090 2.4230 ;
      RECT 0.3310 2.2130 0.7090 2.2630 ;
      RECT 0.6590 2.1630 0.7090 2.2130 ;
      RECT 0.8870 2.0370 0.9370 2.1130 ;
      RECT 0.7350 2.4730 0.7850 2.6900 ;
      RECT 0.6590 2.1130 0.9370 2.1630 ;
      RECT 1.6470 1.2550 1.6970 1.5640 ;
      RECT 1.5710 1.2050 1.6970 1.2550 ;
      RECT 1.5710 1.0620 1.6210 1.2050 ;
      RECT 1.2510 1.9430 1.8070 1.9930 ;
      RECT 0.4740 1.7650 1.6370 1.8150 ;
      RECT 1.0390 1.8150 1.0890 2.0630 ;
      RECT 1.0390 1.7520 1.0890 1.7650 ;
      RECT 0.7350 1.8150 0.7850 2.0630 ;
    LAYER PO ;
      RECT 0.2130 0.0890 0.2430 2.7800 ;
      RECT 1.2770 0.0680 1.3070 2.7800 ;
      RECT 2.1890 0.0670 2.2190 2.7800 ;
      RECT 1.8850 0.0670 1.9150 2.7800 ;
      RECT 2.0370 0.0670 2.0670 2.7800 ;
      RECT 1.4290 0.0680 1.4590 2.7960 ;
      RECT 1.7330 0.0670 1.7630 2.7800 ;
      RECT 1.5810 0.0590 1.6110 2.7800 ;
      RECT 0.3650 0.9880 0.3950 2.7800 ;
      RECT 0.8210 0.0860 0.8510 1.7120 ;
      RECT 1.1250 0.0680 1.1550 2.7780 ;
      RECT 0.6690 0.0890 0.6990 0.7890 ;
      RECT 0.8210 1.8120 0.8510 2.9270 ;
      RECT 0.9730 0.0680 1.0030 1.6680 ;
      RECT 0.3650 0.0870 0.3950 0.8880 ;
      RECT 0.9730 1.7690 1.0030 2.7820 ;
      RECT 0.6690 0.9880 0.6990 2.9300 ;
      RECT 0.5170 0.0780 0.5470 2.7800 ;
      RECT 0.0610 0.0890 0.0910 2.7800 ;
  END
END LSUPENX1_LVT

MACRO LSUPENX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.04 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7940 2.2130 1.1600 2.2630 ;
        RECT 0.9970 2.2630 1.1600 2.3650 ;
    END
    ANTENNAGATEAREA 0.0534 ;
  END A

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.0400 1.7020 ;
        RECT 2.6820 1.7020 2.7920 1.7760 ;
        RECT 2.6820 1.5690 2.7920 1.6420 ;
        RECT 1.0390 1.3520 1.0890 1.6420 ;
        RECT 1.4950 1.4630 1.5450 1.6420 ;
        RECT 2.7110 1.3030 2.7610 1.5690 ;
    END
  END VSS

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 3.0100 3.0400 3.0700 ;
        RECT 1.9220 3.0700 2.0320 3.1440 ;
        RECT 1.9220 2.9370 2.0320 3.0100 ;
        RECT 1.1910 2.5200 1.2410 3.0100 ;
        RECT 0.9110 2.7350 0.9610 3.0100 ;
        RECT 0.8870 2.6740 0.9610 2.7350 ;
        RECT 0.8870 2.5250 0.9370 2.6740 ;
    END
  END VDDL

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3130 2.2240 1.4950 2.3350 ;
    END
    ANTENNAGATEAREA 0.0249 ;
  END EN

  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.0400 0.0300 ;
        RECT 0.4310 0.0300 0.4810 0.4640 ;
        RECT 0.5830 0.0300 0.6330 0.4590 ;
        RECT 1.0390 0.0300 1.0890 0.7210 ;
        RECT 1.9510 0.0300 2.0010 0.9370 ;
        RECT 2.7110 0.0300 2.7610 0.5260 ;
        RECT 2.4070 0.0300 2.4570 0.6610 ;
        RECT 1.7990 0.0300 1.8490 0.2710 ;
        RECT 1.4950 0.2710 1.8490 0.3210 ;
        RECT 1.4950 0.3210 1.5450 0.9050 ;
        RECT 1.7990 0.3210 1.8490 0.9100 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 3.0400 3.3740 ;
    END
  END VDDH

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6190 1.0090 2.7910 1.0590 ;
        RECT 2.6790 1.0590 2.7910 1.1190 ;
        RECT 2.6790 0.8450 2.7290 1.0090 ;
        RECT 2.6790 1.1190 2.7290 1.1780 ;
        RECT 2.2550 0.7950 2.7290 0.8450 ;
        RECT 2.2550 1.1780 2.7290 1.2280 ;
        RECT 2.5590 0.1190 2.6090 0.7950 ;
        RECT 2.2550 0.1190 2.3050 0.7950 ;
        RECT 2.2550 1.2280 2.3050 1.4440 ;
        RECT 2.5590 1.2280 2.6090 1.4440 ;
    END
    ANTENNADIFFAREA 0.412 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1150 -0.1150 3.1550 0.9930 ;
      RECT -0.1150 3.2240 3.1550 3.4590 ;
      RECT -0.1150 2.3510 0.1150 3.2240 ;
      RECT 2.9250 2.3510 3.1550 3.2240 ;
      RECT 0.5750 2.2340 1.4250 2.7640 ;
    LAYER M1 ;
      RECT 0.2390 0.6920 0.7250 0.7420 ;
      RECT 0.2390 0.6840 0.3290 0.6920 ;
      RECT 0.2390 0.7420 0.2890 0.9730 ;
      RECT 0.2790 0.2800 0.3290 0.6840 ;
      RECT 0.2390 0.9730 0.3290 1.0970 ;
      RECT 0.2790 1.0970 0.3290 1.5080 ;
      RECT 1.1930 0.1140 1.6370 0.1280 ;
      RECT 1.1910 0.1280 1.6370 0.1640 ;
      RECT 0.8870 0.1140 0.9370 0.8690 ;
      RECT 1.1910 0.1640 1.2410 0.8690 ;
      RECT 0.8870 0.8690 1.2410 0.9190 ;
      RECT 0.7350 1.0240 1.3330 1.0510 ;
      RECT 0.7750 1.0010 1.3330 1.0240 ;
      RECT 0.7350 1.0510 0.8250 1.0970 ;
      RECT 0.7750 0.8690 0.8250 1.0010 ;
      RECT 0.7350 1.0970 0.7850 1.4110 ;
      RECT 0.3390 0.8190 0.8250 0.8690 ;
      RECT 0.7750 0.5510 0.8250 0.8190 ;
      RECT 0.7350 0.5010 0.8250 0.5510 ;
      RECT 0.7350 0.2740 0.7850 0.5010 ;
      RECT 2.1450 1.0780 2.5490 1.1280 ;
      RECT 2.1450 1.1280 2.1950 1.1450 ;
      RECT 2.1450 0.9430 2.1950 1.0780 ;
      RECT 2.1030 1.1450 2.1950 1.1950 ;
      RECT 2.1020 0.8930 2.1950 0.9430 ;
      RECT 2.1030 1.1950 2.1530 1.4720 ;
      RECT 2.1030 0.1170 2.1530 0.8930 ;
      RECT 0.8110 2.8400 0.8610 2.8620 ;
      RECT 0.6420 2.8620 0.8610 2.9120 ;
      RECT 0.8110 2.9120 0.8610 2.9280 ;
      RECT 1.3430 0.8550 1.4330 0.9050 ;
      RECT 1.3430 0.2710 1.3930 0.8550 ;
      RECT 1.3830 0.9050 1.4330 1.1020 ;
      RECT 0.9360 1.1020 1.4330 1.1520 ;
      RECT 1.3430 1.1520 1.3930 1.5690 ;
      RECT 1.1910 1.3000 1.2410 1.5870 ;
      RECT 0.8870 1.2500 1.2410 1.3000 ;
      RECT 0.8870 1.3000 0.9370 1.5250 ;
      RECT 0.4310 1.5250 0.9370 1.5750 ;
      RECT 0.8870 1.5750 0.9370 1.5870 ;
      RECT 0.5830 1.1380 0.6330 1.5250 ;
      RECT 0.4310 1.0010 0.4810 1.5250 ;
      RECT 0.4310 0.9520 0.5730 1.0010 ;
      RECT 0.4340 0.9510 0.5730 0.9520 ;
      RECT 1.0390 2.4730 1.0890 2.6900 ;
      RECT 0.6590 2.4230 1.0890 2.4730 ;
      RECT 0.8870 2.0370 0.9370 2.1130 ;
      RECT 0.6590 2.1130 0.9370 2.1630 ;
      RECT 0.6590 2.2630 0.7090 2.4230 ;
      RECT 0.3310 2.2130 0.7090 2.2630 ;
      RECT 0.6590 2.1630 0.7090 2.2130 ;
      RECT 0.7350 2.4730 0.7850 2.6900 ;
      RECT 0.4740 1.7680 1.9410 1.8180 ;
      RECT 1.0390 1.8180 1.0890 2.0630 ;
      RECT 0.7350 1.8180 0.7850 2.0630 ;
      RECT 1.6470 0.9940 2.0930 1.0440 ;
      RECT 1.6470 1.0440 1.6970 1.5750 ;
      RECT 1.6470 0.8150 1.6970 0.9940 ;
      RECT 1.2510 1.9430 1.8070 1.9930 ;
      RECT 2.4070 1.4100 2.4570 1.5410 ;
      RECT 1.7980 1.5410 2.4570 1.5840 ;
      RECT 1.7980 1.5840 2.4560 1.5910 ;
      RECT 1.7990 1.1440 1.8490 1.5410 ;
      RECT 1.9510 1.3210 2.0010 1.5410 ;
      RECT 1.7990 1.0940 1.9410 1.1440 ;
      RECT 1.5550 2.0970 2.7010 2.1470 ;
    LAYER PO ;
      RECT 2.9490 0.0670 2.9790 2.7800 ;
      RECT 1.2770 0.0680 1.3070 2.7800 ;
      RECT 0.2130 0.0890 0.2430 2.7800 ;
      RECT 0.5170 0.0780 0.5470 2.7800 ;
      RECT 0.0610 0.0890 0.0910 2.7800 ;
      RECT 0.6690 0.9880 0.6990 2.9300 ;
      RECT 0.9730 1.7690 1.0030 2.7820 ;
      RECT 0.3650 0.0870 0.3950 0.8880 ;
      RECT 0.9730 0.0680 1.0030 1.6680 ;
      RECT 0.8210 1.8120 0.8510 2.9270 ;
      RECT 0.6690 0.0890 0.6990 0.7890 ;
      RECT 1.1250 0.0680 1.1550 2.7780 ;
      RECT 0.8210 0.0860 0.8510 1.7120 ;
      RECT 1.8850 0.0890 1.9150 2.7800 ;
      RECT 0.3650 0.9880 0.3950 2.7800 ;
      RECT 2.0370 0.0670 2.0670 2.7800 ;
      RECT 1.5810 0.0590 1.6110 2.7800 ;
      RECT 1.7330 0.0740 1.7630 2.7800 ;
      RECT 2.1890 0.0670 2.2190 2.7800 ;
      RECT 2.3410 0.0670 2.3710 2.7800 ;
      RECT 2.4930 0.0670 2.5230 2.7800 ;
      RECT 1.4290 0.0680 1.4590 2.7960 ;
      RECT 2.7970 0.0670 2.8270 2.7800 ;
      RECT 2.6450 0.0670 2.6750 2.7800 ;
  END
END LSUPENX2_LVT

MACRO LSUPENX4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.648 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2270 1.0090 3.3990 1.0590 ;
        RECT 3.2870 1.0590 3.3990 1.1190 ;
        RECT 3.2870 0.8450 3.3370 1.0090 ;
        RECT 3.2870 1.1190 3.3370 1.1780 ;
        RECT 2.5590 0.7950 3.3370 0.8450 ;
        RECT 2.5590 1.1780 3.3370 1.2280 ;
        RECT 2.5590 0.1190 2.6090 0.7950 ;
        RECT 2.8630 0.1190 2.9130 0.7950 ;
        RECT 3.1670 0.1190 3.2170 0.7950 ;
        RECT 3.1670 1.2280 3.2170 1.3520 ;
        RECT 2.8630 1.2280 2.9130 1.3520 ;
        RECT 2.5590 1.2280 2.6090 1.3520 ;
    END
    ANTENNADIFFAREA 0.6584 ;
  END Y

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6170 2.2250 1.7990 2.3350 ;
    END
    ANTENNAGATEAREA 0.0255 ;
  END EN

  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.6480 0.0300 ;
        RECT 1.3430 0.0300 1.3930 0.7220 ;
        RECT 2.2550 0.0300 2.3050 0.9370 ;
        RECT 1.0390 0.0300 1.0890 0.7210 ;
        RECT 0.5830 0.0300 0.6330 0.4590 ;
        RECT 0.4310 0.0300 0.4810 0.4640 ;
        RECT 2.7110 0.0300 2.7610 0.6610 ;
        RECT 3.0150 0.0300 3.0650 0.6610 ;
        RECT 3.3190 0.0300 3.3690 0.5260 ;
        RECT 2.1030 0.0300 2.1530 0.2710 ;
        RECT 1.7990 0.2710 2.1530 0.3210 ;
        RECT 1.7990 0.3210 1.8490 0.9050 ;
        RECT 2.1030 0.3210 2.1530 0.9100 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 3.6480 3.3740 ;
    END
  END VDDH

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 3.0100 3.6480 3.0700 ;
        RECT 2.3780 3.0700 2.4880 3.1440 ;
        RECT 2.3780 2.9370 2.4880 3.0100 ;
        RECT 1.1910 2.5200 1.2410 3.0100 ;
        RECT 0.9110 2.7350 0.9610 3.0100 ;
        RECT 0.8870 2.6740 0.9610 2.7350 ;
        RECT 0.8870 2.5250 0.9370 2.6740 ;
    END
  END VDDL

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.6480 1.7020 ;
        RECT 3.2900 1.7020 3.4000 1.7760 ;
        RECT 3.2900 1.5690 3.4000 1.6420 ;
        RECT 1.7990 1.4700 1.8490 1.6420 ;
        RECT 1.3430 1.3520 1.3930 1.6420 ;
        RECT 1.0390 1.3520 1.0890 1.6420 ;
        RECT 3.3190 1.3030 3.3690 1.5690 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7940 2.2130 1.1600 2.2630 ;
        RECT 0.9970 2.2630 1.1600 2.3650 ;
    END
    ANTENNAGATEAREA 0.0501 ;
  END A
  OBS
    LAYER NWELL ;
      RECT -0.1150 3.2240 3.7630 3.4590 ;
      RECT -0.1150 2.3510 0.1150 3.2240 ;
      RECT 3.5330 2.3510 3.7630 3.2240 ;
      RECT 0.5750 2.2340 1.4250 2.7640 ;
      RECT -0.1150 -0.1150 3.7630 0.9930 ;
    LAYER M1 ;
      RECT 0.9360 1.1020 1.7370 1.1520 ;
      RECT 1.6470 1.1520 1.6970 1.5820 ;
      RECT 1.6870 0.9050 1.7370 1.1020 ;
      RECT 1.6470 0.8550 1.7370 0.9050 ;
      RECT 1.6470 0.2710 1.6970 0.8550 ;
      RECT 1.4950 0.1140 1.9410 0.1640 ;
      RECT 0.8870 0.1140 0.9370 0.8690 ;
      RECT 1.1910 0.1280 1.2410 0.8690 ;
      RECT 1.4950 0.1640 1.5450 0.8690 ;
      RECT 0.8870 0.8690 1.5450 0.9190 ;
      RECT 0.8110 2.8400 0.8610 2.8620 ;
      RECT 0.6420 2.8620 0.8610 2.9120 ;
      RECT 0.8110 2.9120 0.8610 2.9280 ;
      RECT 2.4490 1.0780 3.1570 1.1280 ;
      RECT 2.4490 0.9430 2.4990 1.0780 ;
      RECT 2.4490 1.1280 2.4990 1.1450 ;
      RECT 2.4060 0.8930 2.4990 0.9430 ;
      RECT 2.4070 1.1450 2.4990 1.1950 ;
      RECT 2.4070 0.1170 2.4570 0.8930 ;
      RECT 2.4070 1.1950 2.4570 1.3740 ;
      RECT 0.7350 1.0140 1.6370 1.0510 ;
      RECT 0.7750 1.0010 1.6370 1.0140 ;
      RECT 0.7350 1.0510 0.8250 1.0870 ;
      RECT 0.7750 0.9120 0.8250 1.0010 ;
      RECT 0.7350 1.0870 0.7850 1.3900 ;
      RECT 0.3390 0.8620 0.8250 0.9120 ;
      RECT 0.7750 0.5510 0.8250 0.8620 ;
      RECT 0.7350 0.5010 0.8250 0.5510 ;
      RECT 0.7350 0.2740 0.7850 0.5010 ;
      RECT 0.2390 0.6920 0.7250 0.7420 ;
      RECT 0.2390 0.7420 0.2890 1.2240 ;
      RECT 0.2390 0.6840 0.3290 0.6920 ;
      RECT 0.2390 1.2240 0.3290 1.2740 ;
      RECT 0.2790 0.2800 0.3290 0.6840 ;
      RECT 0.2790 1.2740 0.3290 1.5820 ;
      RECT 1.8590 2.0970 3.3090 2.1470 ;
      RECT 0.8870 1.2500 1.5450 1.3000 ;
      RECT 1.4950 1.3000 1.5450 1.5690 ;
      RECT 0.8870 1.3000 0.9370 1.5180 ;
      RECT 0.4310 1.5180 0.9370 1.5670 ;
      RECT 0.5830 1.3230 0.6330 1.5180 ;
      RECT 0.4520 1.5670 0.9370 1.5680 ;
      RECT 0.4310 1.1140 0.4810 1.5180 ;
      RECT 0.4310 1.0640 0.5730 1.1140 ;
      RECT 1.1910 1.3000 1.2410 1.5730 ;
      RECT 0.4740 1.7870 2.2450 1.8370 ;
      RECT 0.7350 1.8370 0.7850 2.0630 ;
      RECT 0.7350 1.7520 0.7850 1.7870 ;
      RECT 1.0390 1.8370 1.0890 2.0760 ;
      RECT 2.1030 1.4240 3.2410 1.4740 ;
      RECT 2.2550 1.4740 2.3050 1.5790 ;
      RECT 2.2550 1.4050 2.3050 1.4240 ;
      RECT 2.1030 1.4740 2.1530 1.5830 ;
      RECT 2.1030 1.1440 2.1530 1.4240 ;
      RECT 2.1030 1.0940 2.2450 1.1440 ;
      RECT 2.7110 1.4740 2.7610 1.5820 ;
      RECT 2.7110 1.4080 2.7610 1.4240 ;
      RECT 3.0150 1.4740 3.0650 1.5780 ;
      RECT 3.0150 1.4040 3.0650 1.4240 ;
      RECT 0.6590 2.4230 1.0890 2.4730 ;
      RECT 1.0390 2.4730 1.0890 2.6900 ;
      RECT 0.6590 2.2630 0.7090 2.4230 ;
      RECT 0.3310 2.2130 0.7090 2.2630 ;
      RECT 0.6590 2.1630 0.7090 2.2130 ;
      RECT 0.8870 2.0370 0.9370 2.1130 ;
      RECT 0.7350 2.4730 0.7850 2.6900 ;
      RECT 0.6590 2.1130 0.9370 2.1630 ;
      RECT 1.9510 0.9940 2.3970 1.0440 ;
      RECT 1.9510 1.0440 2.0010 1.5760 ;
      RECT 1.9510 0.7260 2.0010 0.9940 ;
      RECT 1.5550 1.9430 2.1110 1.9930 ;
    LAYER PO ;
      RECT 2.4930 0.0670 2.5230 2.7800 ;
      RECT 2.0370 0.0740 2.0670 2.7800 ;
      RECT 1.8850 0.0590 1.9150 2.7800 ;
      RECT 2.3410 0.0670 2.3710 2.7800 ;
      RECT 0.3650 1.0980 0.3950 2.7800 ;
      RECT 2.1890 0.0890 2.2190 2.7800 ;
      RECT 0.8210 0.0860 0.8510 1.7120 ;
      RECT 1.1250 0.0680 1.1550 2.7780 ;
      RECT 0.6690 0.0890 0.6990 0.9980 ;
      RECT 0.8210 1.8120 0.8510 2.9270 ;
      RECT 0.9730 0.0680 1.0030 1.6680 ;
      RECT 1.2770 0.0680 1.3070 2.7800 ;
      RECT 1.4290 0.0680 1.4590 2.7800 ;
      RECT 0.3650 0.0870 0.3950 0.9600 ;
      RECT 0.9730 1.7690 1.0030 2.7820 ;
      RECT 0.6690 1.0980 0.6990 2.9300 ;
      RECT 0.5170 0.0780 0.5470 2.7800 ;
      RECT 0.2130 0.0890 0.2430 2.7800 ;
      RECT 0.0610 0.0890 0.0910 2.7800 ;
      RECT 1.5810 0.0680 1.6110 2.7800 ;
      RECT 3.5570 0.0670 3.5870 2.7800 ;
      RECT 3.2530 0.0670 3.2830 2.7800 ;
      RECT 3.4050 0.0670 3.4350 2.7800 ;
      RECT 1.7330 0.0680 1.7630 2.7960 ;
      RECT 2.9490 0.0670 2.9790 2.7800 ;
      RECT 3.1010 0.0670 3.1310 2.7800 ;
      RECT 2.7970 0.0670 2.8270 2.7800 ;
      RECT 2.6450 0.0670 2.6750 2.7800 ;
  END
END LSUPENX4_LVT

MACRO LSUPENX8_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.016 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7940 2.2130 1.1600 2.2630 ;
        RECT 0.9970 2.2630 1.1600 2.3650 ;
    END
    ANTENNAGATEAREA 0.0492 ;
  END A

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 5.0160 1.7020 ;
        RECT 4.6580 1.7020 4.7680 1.7760 ;
        RECT 4.6580 1.5690 4.7680 1.6420 ;
        RECT 1.0390 1.3520 1.0890 1.6420 ;
        RECT 1.9510 1.3520 2.0010 1.6420 ;
        RECT 1.3430 1.3520 1.3930 1.6420 ;
        RECT 1.6470 1.3520 1.6970 1.6420 ;
        RECT 2.4070 1.3420 2.4570 1.6420 ;
        RECT 4.6870 1.3030 4.7370 1.5690 ;
    END
  END VSS

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 3.0100 5.0160 3.0700 ;
        RECT 2.6820 3.0700 2.7920 3.1440 ;
        RECT 2.6820 2.9370 2.7920 3.0100 ;
        RECT 1.1910 2.5200 1.2410 3.0100 ;
        RECT 0.9110 2.7350 0.9610 3.0100 ;
        RECT 0.8870 2.6740 0.9610 2.7350 ;
        RECT 0.8870 2.5250 0.9370 2.6740 ;
    END
  END VDDL

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2250 2.2250 2.4070 2.3350 ;
    END
    ANTENNAGATEAREA 0.027 ;
  END EN

  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 5.0160 0.0300 ;
        RECT 0.4310 0.0300 0.4810 0.4640 ;
        RECT 0.5830 0.0300 0.6330 0.4590 ;
        RECT 1.0390 0.0300 1.0890 0.7210 ;
        RECT 3.0150 0.0300 3.0650 0.8430 ;
        RECT 3.4710 0.0300 3.5210 0.7530 ;
        RECT 4.3830 0.0300 4.4330 0.7530 ;
        RECT 4.0790 0.0300 4.1290 0.7530 ;
        RECT 3.7750 0.0300 3.8250 0.7530 ;
        RECT 1.3430 0.0300 1.3930 0.7220 ;
        RECT 1.6470 0.0300 1.6970 0.7210 ;
        RECT 1.9510 0.0300 2.0010 0.7210 ;
        RECT 4.6880 0.0300 4.7380 0.5260 ;
        RECT 2.7110 0.0300 2.7610 0.2710 ;
        RECT 2.4070 0.2710 2.7610 0.3210 ;
        RECT 2.4070 0.3210 2.4570 0.9050 ;
        RECT 2.7110 0.3210 2.7610 0.9100 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 5.0160 3.3740 ;
    END
  END VDDH

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.5590 0.9370 4.6090 1.0090 ;
        RECT 4.5590 1.0090 4.7670 1.1190 ;
        RECT 3.3190 0.8870 4.6090 0.9370 ;
        RECT 4.5590 1.1190 4.6090 1.1780 ;
        RECT 4.5350 0.1190 4.5850 0.8870 ;
        RECT 4.2310 0.1190 4.2810 0.8870 ;
        RECT 3.6230 0.1190 3.6730 0.8870 ;
        RECT 3.3190 0.1190 3.3690 0.8870 ;
        RECT 3.9270 0.1190 3.9770 0.8870 ;
        RECT 3.3190 1.1780 4.6090 1.2280 ;
        RECT 3.3190 1.2280 3.3690 1.3520 ;
        RECT 3.6230 1.2280 3.6730 1.3520 ;
        RECT 4.2310 1.2280 4.2810 1.3520 ;
        RECT 3.9270 1.2280 3.9770 1.3520 ;
        RECT 4.5350 1.2280 4.6090 1.2600 ;
        RECT 4.5350 1.2600 4.5850 1.3520 ;
    END
    ANTENNADIFFAREA 1.1512 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1150 -0.1150 5.1310 0.9930 ;
      RECT -0.1150 3.2240 5.1310 3.4590 ;
      RECT 4.9010 2.3510 5.1310 3.2240 ;
      RECT -0.1150 2.3510 0.1150 3.2240 ;
      RECT 0.5750 2.2340 1.4250 2.7640 ;
    LAYER M1 ;
      RECT 4.3830 1.4740 4.4330 1.5670 ;
      RECT 2.7110 1.4240 4.4330 1.4740 ;
      RECT 4.3830 1.3930 4.4330 1.4240 ;
      RECT 2.7110 1.4740 2.7610 1.5760 ;
      RECT 3.0150 1.4740 3.0650 1.5720 ;
      RECT 3.0150 1.3980 3.0650 1.4240 ;
      RECT 2.7110 1.1440 2.7610 1.4240 ;
      RECT 2.7110 1.0940 2.8530 1.1440 ;
      RECT 3.4710 1.4740 3.5210 1.5650 ;
      RECT 3.4710 1.3910 3.5210 1.4240 ;
      RECT 3.7750 1.4740 3.8250 1.5660 ;
      RECT 3.7750 1.3920 3.8250 1.4240 ;
      RECT 4.0790 1.4740 4.1290 1.5670 ;
      RECT 4.0790 1.3930 4.1290 1.4240 ;
      RECT 2.1630 1.9430 2.7190 1.9930 ;
      RECT 3.2070 1.0380 4.5090 1.0880 ;
      RECT 4.4590 1.0880 4.5090 1.1230 ;
      RECT 4.4590 0.9980 4.5090 1.0380 ;
      RECT 2.8630 1.2500 2.9130 1.3740 ;
      RECT 2.8630 0.1190 2.9130 0.8940 ;
      RECT 3.2070 1.0880 3.2570 1.2000 ;
      RECT 3.2070 0.9440 3.2570 1.0380 ;
      RECT 2.8630 1.2000 3.2570 1.2500 ;
      RECT 2.8630 0.8940 3.2570 0.9440 ;
      RECT 3.1670 1.2500 3.2170 1.3740 ;
      RECT 3.1670 0.1190 3.2170 0.8940 ;
      RECT 0.2390 0.6920 0.7250 0.7420 ;
      RECT 0.2390 0.6840 0.3290 0.6920 ;
      RECT 0.2390 0.7420 0.2890 1.2230 ;
      RECT 0.2790 0.2800 0.3290 0.6840 ;
      RECT 0.2390 1.2230 0.3290 1.2740 ;
      RECT 0.2790 1.2740 0.3290 1.5810 ;
      RECT 2.1030 0.1140 2.5560 0.1640 ;
      RECT 0.8870 0.1140 0.9370 0.8690 ;
      RECT 1.1910 0.1280 1.2410 0.8690 ;
      RECT 1.4950 0.1280 1.5450 0.8690 ;
      RECT 1.7990 0.1280 1.8490 0.8690 ;
      RECT 2.1030 0.1640 2.1530 0.8690 ;
      RECT 0.8870 0.8690 2.1530 0.9190 ;
      RECT 0.7350 1.0140 2.2450 1.0510 ;
      RECT 0.7750 1.0010 2.2450 1.0140 ;
      RECT 0.7350 1.0510 0.8250 1.0870 ;
      RECT 0.7750 0.9120 0.8250 1.0010 ;
      RECT 0.7350 1.0870 0.7850 1.3900 ;
      RECT 0.3390 0.8620 0.8250 0.9120 ;
      RECT 0.7750 0.5510 0.8250 0.8620 ;
      RECT 0.7350 0.5010 0.8250 0.5510 ;
      RECT 0.7350 0.2740 0.7850 0.5010 ;
      RECT 0.8110 2.8400 0.8610 2.8620 ;
      RECT 0.6420 2.8620 0.8610 2.9120 ;
      RECT 0.8110 2.9120 0.8610 2.9280 ;
      RECT 2.2550 0.8550 2.3450 0.9050 ;
      RECT 2.2550 0.2710 2.3050 0.8550 ;
      RECT 2.2950 0.9050 2.3450 1.1020 ;
      RECT 0.9360 1.1020 2.3450 1.1520 ;
      RECT 2.2550 1.1520 2.3050 1.5660 ;
      RECT 2.1030 1.3000 2.1530 1.5750 ;
      RECT 0.8870 1.2500 2.1530 1.3000 ;
      RECT 0.8870 1.3000 0.9370 1.5090 ;
      RECT 0.4310 1.5090 0.9370 1.5580 ;
      RECT 0.5830 1.3250 0.6330 1.5090 ;
      RECT 0.4520 1.5580 0.9370 1.5590 ;
      RECT 0.4310 1.1300 0.4810 1.5090 ;
      RECT 0.5830 1.5590 0.6330 1.5640 ;
      RECT 0.4310 1.0800 0.5730 1.1300 ;
      RECT 1.1910 1.3000 1.2410 1.5690 ;
      RECT 1.4950 1.3000 1.5450 1.5760 ;
      RECT 1.7990 1.3000 1.8490 1.5730 ;
      RECT 2.4670 2.0970 4.6770 2.1470 ;
      RECT 1.0390 2.4730 1.0890 2.6900 ;
      RECT 0.6590 2.4230 1.0890 2.4730 ;
      RECT 0.8870 2.0370 0.9370 2.1130 ;
      RECT 0.6590 2.1130 0.9370 2.1630 ;
      RECT 0.6590 2.2630 0.7090 2.4230 ;
      RECT 0.3310 2.2130 0.7090 2.2630 ;
      RECT 0.6590 2.1630 0.7090 2.2130 ;
      RECT 0.7350 2.4730 0.7850 2.6900 ;
      RECT 0.4740 1.7880 2.8530 1.8380 ;
      RECT 1.0390 1.8380 1.0890 2.0630 ;
      RECT 0.7350 1.8380 0.7850 2.0630 ;
      RECT 2.5590 0.9940 3.1570 1.0440 ;
      RECT 2.5590 1.0440 2.6090 1.5710 ;
      RECT 2.5590 0.7370 2.6090 0.9940 ;
    LAYER PO ;
      RECT 0.2130 0.0890 0.2430 2.7800 ;
      RECT 0.5170 0.0780 0.5470 2.7800 ;
      RECT 0.0610 0.0890 0.0910 2.7800 ;
      RECT 0.6690 1.1280 0.6990 2.9300 ;
      RECT 0.9730 1.7690 1.0030 2.7820 ;
      RECT 1.7330 0.0680 1.7630 2.7800 ;
      RECT 0.3650 0.0870 0.3950 0.9600 ;
      RECT 2.0370 0.0680 2.0670 2.7800 ;
      RECT 1.4290 0.0680 1.4590 2.7800 ;
      RECT 1.2770 0.0680 1.3070 2.7800 ;
      RECT 1.5810 0.0680 1.6110 2.7800 ;
      RECT 0.9730 0.0680 1.0030 1.6680 ;
      RECT 0.8210 1.8120 0.8510 2.9270 ;
      RECT 1.8850 0.0680 1.9150 2.7800 ;
      RECT 0.6690 0.0890 0.6990 1.0250 ;
      RECT 1.1250 0.0680 1.1550 2.7780 ;
      RECT 0.8210 0.0860 0.8510 1.7120 ;
      RECT 2.7970 0.0890 2.8270 2.7800 ;
      RECT 0.3650 1.1280 0.3950 2.7800 ;
      RECT 2.9490 0.0670 2.9790 2.7800 ;
      RECT 2.4930 0.0590 2.5230 2.7800 ;
      RECT 2.6450 0.0740 2.6750 2.7800 ;
      RECT 3.2530 0.0670 3.2830 2.7800 ;
      RECT 3.1010 0.0670 3.1310 2.7800 ;
      RECT 3.4050 0.0670 3.4350 2.7800 ;
      RECT 3.5570 0.0670 3.5870 2.7800 ;
      RECT 3.8610 0.0670 3.8910 2.7800 ;
      RECT 3.7090 0.0670 3.7390 2.7800 ;
      RECT 4.1650 0.0670 4.1950 2.7800 ;
      RECT 4.0130 0.0670 4.0430 2.7800 ;
      RECT 4.3170 0.0670 4.3470 2.7800 ;
      RECT 4.4690 0.0670 4.4990 2.7800 ;
      RECT 2.3410 0.0680 2.3710 2.7960 ;
      RECT 4.7730 0.0670 4.8030 2.7800 ;
      RECT 4.6210 0.0670 4.6510 2.7800 ;
      RECT 4.9250 0.0670 4.9550 2.7800 ;
      RECT 2.1890 0.0680 2.2190 2.7800 ;
  END
END LSUPENX8_LVT

MACRO LSDNENCLX4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.584 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.5840 0.0300 ;
        RECT 1.6470 0.0300 1.6970 0.3450 ;
        RECT 1.9510 0.0300 2.0010 0.3450 ;
        RECT 1.3430 0.0300 1.3930 0.3450 ;
        RECT 0.8870 0.0300 0.9370 0.5050 ;
        RECT 2.2550 0.0300 2.3050 0.4850 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 2.5840 3.3740 ;
    END
  END VDDL

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7900 1.1470 0.9810 1.2810 ;
    END
    ANTENNAGATEAREA 0.063 ;
  END EN

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.5840 1.7020 ;
        RECT 0.0980 1.7020 0.2080 1.7750 ;
        RECT 0.0980 1.5680 0.2080 1.6420 ;
        RECT 0.4310 1.4960 0.4810 1.6420 ;
        RECT 1.6470 1.3630 1.6970 1.6420 ;
        RECT 1.9510 1.3630 2.0010 1.6420 ;
        RECT 1.3430 1.5220 1.3930 1.6420 ;
        RECT 2.2550 1.3270 2.3050 1.6420 ;
        RECT 1.0390 1.7020 1.0890 2.1290 ;
        RECT 0.8870 1.5170 0.9370 1.6420 ;
    END
  END VSS

  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 3.0100 2.5840 3.0700 ;
        RECT 1.3140 3.0700 1.4240 3.1430 ;
        RECT 1.3140 2.9360 1.4240 3.0100 ;
        RECT 1.0390 2.5250 1.0890 3.0100 ;
        RECT 1.3430 2.5200 1.3930 2.9360 ;
    END
  END VDDH

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.1710 0.6700 2.2210 0.6940 ;
        RECT 2.1710 0.6940 2.3630 0.8280 ;
        RECT 1.4950 0.6200 2.2210 0.6700 ;
        RECT 2.1710 0.8280 2.2210 1.1610 ;
        RECT 2.1030 0.2170 2.1530 0.6200 ;
        RECT 1.4950 0.1850 1.5450 0.6200 ;
        RECT 1.7990 0.2170 1.8490 0.6200 ;
        RECT 1.4950 1.1610 2.2210 1.2110 ;
        RECT 2.1030 1.2110 2.1530 1.5830 ;
        RECT 1.4950 1.2110 1.5450 1.5830 ;
        RECT 1.7990 1.2110 1.8490 1.5830 ;
    END
    ANTENNADIFFAREA 0.3976 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9460 2.2130 1.3120 2.2630 ;
        RECT 1.1490 2.2630 1.3120 2.3650 ;
    END
    ANTENNAGATEAREA 0.0261 ;
  END A
  OBS
    LAYER NWELL ;
      RECT 0.5750 2.2340 1.6170 2.7640 ;
      RECT -0.1150 3.2240 2.6990 3.4590 ;
      RECT -0.1150 2.3510 0.1150 3.2240 ;
      RECT 2.4690 2.3510 2.6990 3.2240 ;
      RECT -0.1150 -0.1150 2.6990 0.9930 ;
    LAYER M1 ;
      RECT 0.7350 0.6640 1.0890 0.7140 ;
      RECT 1.0390 0.2300 1.0890 0.6640 ;
      RECT 0.7350 0.1380 0.7850 0.6640 ;
      RECT 0.4310 0.0880 0.7850 0.1380 ;
      RECT 0.4310 0.1380 0.4810 0.6310 ;
      RECT 1.3830 1.0330 2.0930 1.0830 ;
      RECT 1.3830 1.0830 1.4330 1.2010 ;
      RECT 1.3830 0.8510 1.4330 1.0330 ;
      RECT 1.1910 1.2010 1.4330 1.2510 ;
      RECT 1.1720 0.8010 1.4330 0.8510 ;
      RECT 1.1910 1.2510 1.2410 1.2950 ;
      RECT 1.2200 1.0280 1.3330 1.0780 ;
      RECT 0.2790 0.2280 0.3290 0.7810 ;
      RECT 0.7350 1.4340 0.7850 1.5840 ;
      RECT 0.6330 0.8310 0.6830 0.9010 ;
      RECT 0.6330 0.9510 0.6830 1.1980 ;
      RECT 0.2790 0.7810 0.6830 0.8310 ;
      RECT 0.5830 1.1980 0.6830 1.2620 ;
      RECT 0.5830 0.2300 0.6330 0.7810 ;
      RECT 0.5830 1.2620 0.6330 1.3840 ;
      RECT 0.5830 1.4340 0.6330 1.5840 ;
      RECT 0.6330 0.9010 1.2700 0.9510 ;
      RECT 1.2200 0.9510 1.2700 1.0280 ;
      RECT 0.5830 1.3840 1.0890 1.4340 ;
      RECT 1.0390 1.4340 1.0890 1.5840 ;
      RECT 0.8270 2.4230 1.2410 2.4730 ;
      RECT 1.1910 2.4730 1.2410 2.6900 ;
      RECT 0.8270 2.2850 0.8770 2.4230 ;
      RECT 0.7660 2.2630 0.8770 2.2850 ;
      RECT 0.3380 2.2130 0.8770 2.2630 ;
      RECT 0.7660 2.1840 0.8770 2.2130 ;
      RECT 0.8270 2.1280 0.8770 2.1840 ;
      RECT 0.8870 2.4730 0.9370 2.6900 ;
      RECT 0.8270 2.0780 0.9370 2.1280 ;
      RECT 0.8870 1.9760 0.9370 2.0780 ;
      RECT 0.7950 1.0280 1.0290 1.0780 ;
      RECT 0.3390 1.0280 0.5730 1.0780 ;
    LAYER PO ;
      RECT 0.6690 0.0780 0.6990 2.7810 ;
      RECT 2.0370 0.0620 2.0670 2.7800 ;
      RECT 2.1890 0.0620 2.2190 2.7800 ;
      RECT 0.3650 0.0890 0.3950 2.7800 ;
      RECT 1.1250 0.0870 1.1550 2.7780 ;
      RECT 2.3410 0.0620 2.3710 2.7800 ;
      RECT 1.8850 0.0620 1.9150 2.7800 ;
      RECT 0.8210 0.0780 0.8510 2.7800 ;
      RECT 1.5810 0.0620 1.6110 2.7800 ;
      RECT 1.2770 0.0680 1.3070 2.7800 ;
      RECT 1.4290 0.0680 1.4590 2.7800 ;
      RECT 2.4930 0.0670 2.5230 2.7800 ;
      RECT 1.7330 0.0620 1.7630 2.7800 ;
      RECT 0.9730 0.0780 1.0030 1.7850 ;
      RECT 0.9730 1.9210 1.0030 2.7820 ;
      RECT 0.2130 0.0890 0.2430 2.7800 ;
      RECT 0.0610 0.0890 0.0910 2.7800 ;
      RECT 0.5170 0.0890 0.5470 2.7800 ;
  END
END LSDNENCLX4_LVT

MACRO LSDNENCLX8_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.344 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.3440 0.0300 ;
        RECT 2.7110 0.0300 2.7610 0.3450 ;
        RECT 1.7990 0.0300 1.8490 0.3450 ;
        RECT 2.4070 0.0300 2.4570 0.3500 ;
        RECT 2.1030 0.0300 2.1530 0.3450 ;
        RECT 1.1910 0.0300 1.2410 0.3450 ;
        RECT 1.4950 0.0300 1.5450 0.3450 ;
        RECT 0.8870 0.0300 0.9370 0.5050 ;
        RECT 3.0150 0.0300 3.0650 0.4850 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 3.3440 3.3740 ;
    END
  END VDDL

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7900 1.0890 0.9810 1.2710 ;
    END
    ANTENNAGATEAREA 0.066 ;
  END EN

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.3440 1.7020 ;
        RECT 2.9860 1.7020 3.0960 1.7750 ;
        RECT 2.9860 1.5680 3.0960 1.6420 ;
        RECT 1.0390 1.7020 1.0890 2.1290 ;
        RECT 0.8870 1.5170 0.9370 1.6420 ;
        RECT 2.7110 1.3630 2.7610 1.6420 ;
        RECT 1.7990 1.3630 1.8490 1.6420 ;
        RECT 2.4070 1.3630 2.4570 1.6420 ;
        RECT 2.1030 1.3630 2.1530 1.6420 ;
        RECT 0.4310 1.5060 0.4810 1.6420 ;
        RECT 1.1910 1.5220 1.2410 1.6420 ;
        RECT 1.4950 1.5260 1.5450 1.6420 ;
        RECT 3.0150 1.3030 3.0650 1.5680 ;
    END
  END VSS

  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 3.0100 3.3440 3.0700 ;
        RECT 1.7700 3.0700 1.8800 3.1430 ;
        RECT 1.7700 2.9360 1.8800 3.0100 ;
        RECT 1.3430 2.5200 1.3930 3.0100 ;
        RECT 1.0390 2.5250 1.0890 3.0100 ;
    END
  END VDDH

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9340 0.6700 2.9840 0.6940 ;
        RECT 2.9340 0.6940 3.1230 0.8280 ;
        RECT 1.6470 0.6200 2.9840 0.6700 ;
        RECT 2.9340 0.8280 2.9840 1.2010 ;
        RECT 2.8630 0.2170 2.9130 0.6200 ;
        RECT 2.2550 0.2170 2.3050 0.6200 ;
        RECT 2.5590 0.1850 2.6090 0.6200 ;
        RECT 1.9510 0.2170 2.0010 0.6200 ;
        RECT 1.6470 0.1850 1.6970 0.6200 ;
        RECT 1.6470 1.2010 2.9840 1.2510 ;
        RECT 2.5590 1.2510 2.6090 1.5730 ;
        RECT 2.8630 1.2510 2.9130 1.5730 ;
        RECT 2.2550 1.2510 2.3050 1.5730 ;
        RECT 1.6470 1.2510 1.6970 1.5730 ;
        RECT 1.9510 1.2510 2.0010 1.5730 ;
    END
    ANTENNADIFFAREA 0.6952 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9460 2.2130 1.3120 2.2630 ;
        RECT 1.1490 2.2630 1.3120 2.3650 ;
    END
    ANTENNAGATEAREA 0.0261 ;
  END A
  OBS
    LAYER NWELL ;
      RECT -0.1150 3.2240 3.4590 3.4580 ;
      RECT -0.1150 2.3510 0.1150 3.2240 ;
      RECT 3.2290 2.3510 3.4590 3.2240 ;
      RECT 0.5750 2.2340 1.6170 2.7640 ;
      RECT -0.1150 -0.1150 3.4590 0.9930 ;
    LAYER M1 ;
      RECT 1.5350 1.0330 2.8840 1.0830 ;
      RECT 1.5350 0.8510 1.5850 1.0330 ;
      RECT 1.5350 1.0830 1.5850 1.2010 ;
      RECT 1.3430 0.8010 1.5850 0.8510 ;
      RECT 1.3430 1.2010 1.5850 1.2510 ;
      RECT 1.3430 0.8510 1.3930 0.9170 ;
      RECT 1.3430 1.2510 1.3930 1.3040 ;
      RECT 1.0390 0.2300 1.0890 0.6640 ;
      RECT 0.7350 0.6640 1.0890 0.7140 ;
      RECT 0.7350 0.1440 0.7850 0.6640 ;
      RECT 0.4310 0.0940 0.7850 0.1440 ;
      RECT 0.4310 0.1440 0.4810 0.6310 ;
      RECT 1.2200 1.0280 1.4850 1.0780 ;
      RECT 0.2790 0.2280 0.3290 0.7810 ;
      RECT 0.7350 1.4330 0.7850 1.5840 ;
      RECT 0.5830 0.2300 0.6330 0.7810 ;
      RECT 0.6330 0.8310 0.6830 1.1980 ;
      RECT 0.5830 1.1980 0.6830 1.2620 ;
      RECT 0.5830 1.2620 0.6330 1.3830 ;
      RECT 0.5830 1.4330 0.6330 1.5840 ;
      RECT 0.5830 1.3830 1.0890 1.4330 ;
      RECT 1.0390 1.4330 1.0890 1.5840 ;
      RECT 1.2200 0.8310 1.2700 1.0280 ;
      RECT 0.2790 0.7810 1.2700 0.8310 ;
      RECT 0.8270 2.4230 1.2410 2.4730 ;
      RECT 1.1910 2.4730 1.2410 2.6900 ;
      RECT 0.8270 2.2850 0.8770 2.4230 ;
      RECT 0.7660 2.2630 0.8770 2.2850 ;
      RECT 0.3380 2.2130 0.8770 2.2630 ;
      RECT 0.7660 2.1840 0.8770 2.2130 ;
      RECT 0.8270 2.1280 0.8770 2.1840 ;
      RECT 0.8870 2.4730 0.9370 2.6900 ;
      RECT 0.8270 2.0780 0.9370 2.1280 ;
      RECT 0.8870 1.9760 0.9370 2.0780 ;
      RECT 0.7950 0.9700 1.0290 1.0200 ;
      RECT 0.3390 1.0280 0.5730 1.0780 ;
    LAYER PO ;
      RECT 3.2530 0.0650 3.2830 2.7800 ;
      RECT 0.6690 0.0780 0.6990 2.7810 ;
      RECT 2.0370 0.0600 2.0670 2.7800 ;
      RECT 2.1890 0.0600 2.2190 2.7800 ;
      RECT 2.3410 0.0600 2.3710 2.7800 ;
      RECT 2.4930 0.0600 2.5230 2.7800 ;
      RECT 2.6450 0.0600 2.6750 2.7800 ;
      RECT 2.7970 0.0600 2.8270 2.7800 ;
      RECT 0.3650 0.0890 0.3950 2.7800 ;
      RECT 1.1250 0.0870 1.1550 2.7780 ;
      RECT 2.9490 0.0600 2.9790 2.7800 ;
      RECT 1.8850 0.0600 1.9150 2.7800 ;
      RECT 0.8210 0.0780 0.8510 2.7800 ;
      RECT 1.5810 0.0600 1.6110 2.7800 ;
      RECT 1.2770 0.0650 1.3070 2.7800 ;
      RECT 1.4290 0.0640 1.4590 2.7800 ;
      RECT 3.1010 0.0650 3.1310 2.7800 ;
      RECT 1.7330 0.0600 1.7630 2.7800 ;
      RECT 0.9730 0.0780 1.0030 1.7850 ;
      RECT 0.9730 1.9210 1.0030 2.7820 ;
      RECT 0.2130 0.0890 0.2430 2.7800 ;
      RECT 0.0610 0.0890 0.0910 2.7800 ;
      RECT 0.5170 0.0890 0.5470 2.7800 ;
  END
END LSDNENCLX8_LVT

MACRO LSDNENSSX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.584 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.1640 0.7060 2.3350 0.8160 ;
    END
    ANTENNAGATEAREA 0.0237 ;
  END EN

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.5840 0.0300 ;
        RECT 2.2550 0.0300 2.3050 0.3690 ;
        RECT 1.6470 0.0300 1.6970 0.3680 ;
        RECT 1.3430 0.0300 1.3930 0.3680 ;
    END
  END VSS

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.5840 1.7020 ;
        RECT 2.2550 1.0780 2.3050 1.6420 ;
        RECT 1.1910 1.2580 1.2410 1.6420 ;
        RECT 0.7350 1.3290 0.7850 1.6420 ;
        RECT 0.4310 1.2190 0.4810 1.6420 ;
    END
  END VDDL

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.8400 0.5110 0.8900 ;
        RECT 0.4010 0.8900 0.5110 0.9670 ;
    END
    ANTENNAGATEAREA 0.0237 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0390 0.8160 1.9030 0.8660 ;
        RECT 1.0390 0.8660 1.0890 1.1090 ;
        RECT 1.3430 0.8660 1.3930 1.2140 ;
        RECT 1.7690 0.8660 1.9030 0.9670 ;
        RECT 1.8530 0.5930 1.9030 0.8160 ;
        RECT 1.0390 0.5430 1.9030 0.5930 ;
        RECT 1.0390 0.1940 1.0890 0.5430 ;
    END
    ANTENNADIFFAREA 0.206 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 2.6990 1.7730 ;
    LAYER M1 ;
      RECT 2.0210 0.5020 2.1530 0.5520 ;
      RECT 2.1030 0.1760 2.1530 0.5020 ;
      RECT 2.0210 0.9100 2.1290 0.9110 ;
      RECT 2.0210 0.9110 2.1530 0.9600 ;
      RECT 2.1030 0.9600 2.1530 1.1650 ;
      RECT 1.6880 1.1650 2.1530 1.2150 ;
      RECT 2.1030 1.2150 2.1530 1.5280 ;
      RECT 2.0210 0.5520 2.0710 0.9100 ;
      RECT 1.1910 0.4400 1.8490 0.4900 ;
      RECT 1.7990 0.1940 1.8490 0.4400 ;
      RECT 1.1910 0.1380 1.2410 0.4400 ;
      RECT 0.4310 0.0880 1.2410 0.1380 ;
      RECT 1.4950 0.1940 1.5450 0.4400 ;
      RECT 0.4310 0.1380 0.4810 0.3690 ;
      RECT 0.7350 0.1380 0.7850 0.3680 ;
      RECT 0.9270 0.6520 1.1810 0.7020 ;
      RECT 0.9270 0.7020 0.9770 0.8040 ;
      RECT 0.9270 0.5820 0.9770 0.6520 ;
      RECT 0.8870 0.8040 0.9770 0.8540 ;
      RECT 0.8870 0.5320 0.9770 0.5820 ;
      RECT 0.8870 0.8540 0.9370 1.0240 ;
      RECT 0.8870 0.1940 0.9370 0.5320 ;
      RECT 0.5830 0.7730 0.8250 0.8230 ;
      RECT 0.5830 0.8230 0.6330 1.2310 ;
      RECT 0.7750 0.7050 0.8250 0.7730 ;
      RECT 0.7750 0.6550 0.8770 0.7050 ;
      RECT 0.7750 0.5510 0.8250 0.6550 ;
      RECT 0.5830 0.5010 0.8250 0.5510 ;
      RECT 0.5830 0.1940 0.6330 0.5010 ;
      RECT 1.2510 0.6530 1.7900 0.7030 ;
      RECT 0.2390 0.6510 0.7250 0.7010 ;
      RECT 0.2790 0.1950 0.3290 0.6510 ;
      RECT 0.2390 0.9470 0.3290 0.9970 ;
      RECT 0.2790 0.9970 0.3290 1.5050 ;
      RECT 0.2390 0.7010 0.2890 0.9470 ;
    LAYER PO ;
      RECT 2.0370 0.1340 2.0670 1.6120 ;
      RECT 1.7330 0.1340 1.7630 1.6120 ;
      RECT 1.8850 0.1330 1.9150 1.6120 ;
      RECT 1.1250 0.1330 1.1550 1.6120 ;
      RECT 1.5810 0.1330 1.6110 1.6120 ;
      RECT 2.4930 0.1330 2.5230 1.6120 ;
      RECT 0.9730 0.1330 1.0030 1.6120 ;
      RECT 1.4290 0.1340 1.4590 1.6120 ;
      RECT 1.2770 0.1340 1.3070 1.6120 ;
      RECT 0.3650 0.1330 0.3950 1.6120 ;
      RECT 0.5170 0.1330 0.5470 1.6120 ;
      RECT 0.8210 0.1330 0.8510 1.6120 ;
      RECT 0.6690 0.1330 0.6990 1.6120 ;
      RECT 0.0610 0.1330 0.0910 1.6040 ;
      RECT 2.1890 0.1340 2.2190 1.6120 ;
      RECT 2.3410 0.1330 2.3710 1.6120 ;
      RECT 0.2130 0.1330 0.2430 1.6120 ;
  END
END LSDNENSSX1_LVT

MACRO LSDNENSSX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.04 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.6290 0.7050 2.7910 0.8260 ;
    END
    ANTENNAGATEAREA 0.0237 ;
  END EN

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.0400 0.0300 ;
        RECT 1.4950 0.0300 1.5450 0.3680 ;
        RECT 1.7990 0.0300 1.8490 0.3680 ;
        RECT 2.7110 0.0300 2.7610 0.4710 ;
        RECT 2.1030 0.0300 2.1530 0.3680 ;
    END
  END VSS

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.0400 1.7020 ;
        RECT 0.4310 1.3170 0.4810 1.6420 ;
        RECT 1.0390 1.3640 1.0890 1.6420 ;
        RECT 0.7350 1.3240 0.7850 1.6420 ;
        RECT 1.3430 1.3360 1.3930 1.6420 ;
        RECT 1.6470 1.0100 1.6970 1.6420 ;
        RECT 2.7110 1.0280 2.7610 1.6420 ;
    END
  END VDDL

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.8360 0.5110 0.8860 ;
        RECT 0.4010 0.8860 0.5110 0.9670 ;
    END
    ANTENNAGATEAREA 0.0237 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1910 0.8660 2.3440 0.8680 ;
        RECT 1.1910 0.8680 1.2410 1.0630 ;
        RECT 1.4950 0.8680 1.5450 1.1100 ;
        RECT 2.2250 0.8680 2.3350 0.9670 ;
        RECT 1.1910 0.8180 2.3770 0.8660 ;
        RECT 2.3270 0.6020 2.3770 0.8180 ;
        RECT 1.1910 0.5520 2.3770 0.6020 ;
        RECT 1.1910 0.1940 1.2410 0.5520 ;
    END
    ANTENNADIFFAREA 0.2464 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 3.1550 1.7730 ;
    LAYER M1 ;
      RECT 0.2390 0.6600 0.7250 0.7100 ;
      RECT 0.2790 0.1950 0.3290 0.6600 ;
      RECT 0.2390 0.9430 0.3290 0.9930 ;
      RECT 0.2790 0.9930 0.3290 1.5010 ;
      RECT 0.2390 0.7100 0.2890 0.9430 ;
      RECT 1.3430 0.4520 2.3050 0.5020 ;
      RECT 2.2550 0.1940 2.3050 0.4520 ;
      RECT 1.3430 0.1380 1.3930 0.4520 ;
      RECT 0.4310 0.0880 1.3930 0.1380 ;
      RECT 1.6470 0.1940 1.6970 0.4520 ;
      RECT 1.9510 0.1940 2.0010 0.4520 ;
      RECT 0.7350 0.1380 0.7850 0.3680 ;
      RECT 1.0390 0.1380 1.0890 0.4600 ;
      RECT 0.4310 0.1380 0.4810 0.4610 ;
      RECT 0.9270 0.6520 1.3330 0.7020 ;
      RECT 0.9270 0.7020 0.9770 0.8040 ;
      RECT 0.9270 0.5820 0.9770 0.6520 ;
      RECT 0.8870 0.8040 0.9770 0.8540 ;
      RECT 0.8870 0.5320 0.9770 0.5820 ;
      RECT 0.8870 0.8540 0.9370 1.0190 ;
      RECT 0.8870 0.1940 0.9370 0.5320 ;
      RECT 0.5830 0.7730 0.8250 0.8230 ;
      RECT 0.5830 0.8230 0.6330 1.0510 ;
      RECT 0.7750 0.7000 0.8250 0.7730 ;
      RECT 0.7750 0.6500 0.8770 0.7000 ;
      RECT 0.7750 0.5510 0.8250 0.6500 ;
      RECT 0.5830 0.5010 0.8250 0.5510 ;
      RECT 0.5830 0.1940 0.6330 0.5010 ;
      RECT 1.4030 0.6530 2.2450 0.7030 ;
      RECT 2.4780 0.9060 2.6070 0.9560 ;
      RECT 2.5570 0.9560 2.6070 1.4450 ;
      RECT 2.1450 1.4450 2.6070 1.4950 ;
      RECT 2.5590 0.1820 2.6090 0.6070 ;
      RECT 2.5570 1.4950 2.6070 1.5250 ;
      RECT 2.4780 0.6070 2.6090 0.6550 ;
      RECT 2.4780 0.6550 2.5790 0.6570 ;
      RECT 2.4780 0.6570 2.5280 0.9060 ;
    LAYER PO ;
      RECT 0.9730 0.1330 1.0030 1.6120 ;
      RECT 0.8210 0.1330 0.8510 1.6120 ;
      RECT 0.6690 0.1330 0.6990 1.6120 ;
      RECT 1.8850 0.1330 1.9150 1.6120 ;
      RECT 2.1890 0.1330 2.2190 1.6120 ;
      RECT 1.7330 0.1340 1.7630 1.6120 ;
      RECT 1.4290 0.1330 1.4590 1.6120 ;
      RECT 1.5810 0.1340 1.6110 1.6120 ;
      RECT 1.1250 0.1330 1.1550 1.6120 ;
      RECT 1.2770 0.1340 1.3070 1.6120 ;
      RECT 0.3650 0.1330 0.3950 1.6120 ;
      RECT 0.5170 0.1330 0.5470 1.6120 ;
      RECT 0.0610 0.1330 0.0910 1.6040 ;
      RECT 0.2130 0.1330 0.2430 1.6120 ;
      RECT 2.6450 0.1330 2.6750 1.6120 ;
      RECT 2.3410 0.1340 2.3710 1.6120 ;
      RECT 2.7970 0.1340 2.8270 1.6120 ;
      RECT 2.0370 0.1340 2.0670 1.6120 ;
      RECT 2.4930 0.1330 2.5230 1.6120 ;
      RECT 2.9490 0.1340 2.9790 1.6120 ;
  END
END LSDNENSSX2_LVT

MACRO LSDNENSSX4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.344 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.3440 0.0300 ;
        RECT 3.0150 0.0300 3.0650 0.4900 ;
        RECT 2.4070 0.0300 2.4570 0.3680 ;
        RECT 2.1030 0.0300 2.1530 0.3680 ;
        RECT 1.7990 0.0300 1.8490 0.3680 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1910 0.8310 2.6980 0.8810 ;
        RECT 2.5290 0.8810 2.6390 0.9680 ;
        RECT 2.1030 0.8810 2.1530 1.2210 ;
        RECT 1.7990 0.8810 1.8490 1.2090 ;
        RECT 1.1910 0.8810 1.2410 1.0540 ;
        RECT 1.4950 0.8810 1.5450 1.0450 ;
        RECT 2.6480 0.5990 2.6980 0.8310 ;
        RECT 1.1910 0.5490 2.6980 0.5990 ;
        RECT 1.1910 0.1940 1.2410 0.5490 ;
        RECT 1.4950 0.1940 1.5450 0.5490 ;
    END
    ANTENNADIFFAREA 0.4928 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.8000 0.5110 0.8500 ;
        RECT 0.4010 0.8500 0.5110 0.9670 ;
    END
    ANTENNAGATEAREA 0.0237 ;
  END A

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9390 0.6430 2.9890 0.6660 ;
        RECT 2.9390 0.6660 3.0950 0.7310 ;
        RECT 2.9850 0.7310 3.0950 0.8150 ;
    END
    ANTENNAGATEAREA 0.0237 ;
  END EN

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.3440 1.7020 ;
        RECT 3.0150 0.9850 3.0650 1.6420 ;
        RECT 1.9510 1.3350 2.0010 1.6420 ;
        RECT 0.4310 1.2790 0.4810 1.6420 ;
        RECT 2.2550 1.0100 2.3050 1.6420 ;
        RECT 0.7350 1.3330 0.7850 1.6420 ;
        RECT 1.0390 1.3150 1.0890 1.6420 ;
        RECT 1.3430 1.3160 1.3930 1.6420 ;
        RECT 1.6470 1.3360 1.6970 1.6420 ;
    END
  END VDDL
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 3.4570 1.7730 ;
    LAYER M1 ;
      RECT 2.8330 0.9640 2.9130 1.0140 ;
      RECT 2.8630 1.0140 2.9130 1.3240 ;
      RECT 2.4490 1.3240 2.9130 1.3740 ;
      RECT 2.8330 0.5300 2.9130 0.5890 ;
      RECT 2.8630 1.3740 2.9130 1.5130 ;
      RECT 2.8630 0.1880 2.9130 0.5300 ;
      RECT 2.8330 0.5890 2.8830 0.9640 ;
      RECT 1.6470 0.4360 2.6090 0.4860 ;
      RECT 2.5590 0.1940 2.6090 0.4360 ;
      RECT 1.6470 0.1380 1.6970 0.4360 ;
      RECT 0.4310 0.0880 1.6970 0.1380 ;
      RECT 1.9510 0.1940 2.0010 0.4360 ;
      RECT 2.2550 0.1940 2.3050 0.4360 ;
      RECT 1.0390 0.1380 1.0890 0.4600 ;
      RECT 0.7350 0.1380 0.7850 0.3680 ;
      RECT 0.4310 0.1380 0.4810 0.4610 ;
      RECT 1.3430 0.1380 1.3930 0.4600 ;
      RECT 0.9270 0.6610 1.6370 0.7110 ;
      RECT 0.9270 0.7110 0.9770 0.8040 ;
      RECT 0.9270 0.5820 0.9770 0.6610 ;
      RECT 0.8870 0.8040 0.9770 0.8540 ;
      RECT 0.8870 0.5320 0.9770 0.5820 ;
      RECT 0.8870 0.8540 0.9370 1.0130 ;
      RECT 0.8870 0.1940 0.9370 0.5320 ;
      RECT 0.2390 0.6600 0.7250 0.7100 ;
      RECT 0.2790 0.1950 0.3290 0.6600 ;
      RECT 0.2390 0.9070 0.3290 0.9570 ;
      RECT 0.2790 0.9570 0.3290 1.4650 ;
      RECT 0.2390 0.7100 0.2890 0.9070 ;
      RECT 0.5830 0.7730 0.8250 0.8230 ;
      RECT 0.5830 0.8230 0.6330 1.0570 ;
      RECT 0.7750 0.7000 0.8250 0.7730 ;
      RECT 0.7750 0.6500 0.8770 0.7000 ;
      RECT 0.7750 0.5510 0.8250 0.6500 ;
      RECT 0.5830 0.5010 0.8250 0.5510 ;
      RECT 0.5830 0.1940 0.6330 0.5010 ;
      RECT 1.7070 0.6600 2.5870 0.7100 ;
    LAYER PO ;
      RECT 0.2130 0.1330 0.2430 1.6120 ;
      RECT 0.0610 0.1330 0.0910 1.6040 ;
      RECT 0.5170 0.1330 0.5470 1.6120 ;
      RECT 0.9730 0.1330 1.0030 1.6120 ;
      RECT 0.3650 0.1330 0.3950 1.6120 ;
      RECT 1.2770 0.1340 1.3070 1.6120 ;
      RECT 1.1250 0.1330 1.1550 1.6120 ;
      RECT 1.5810 0.1340 1.6110 1.6120 ;
      RECT 1.4290 0.1330 1.4590 1.6120 ;
      RECT 1.7330 0.1330 1.7630 1.6120 ;
      RECT 2.0370 0.1340 2.0670 1.6120 ;
      RECT 1.8850 0.1330 1.9150 1.6120 ;
      RECT 2.1890 0.1330 2.2190 1.6120 ;
      RECT 2.3410 0.1330 2.3710 1.6120 ;
      RECT 2.4930 0.1340 2.5230 1.6120 ;
      RECT 0.6690 0.1330 0.6990 1.6120 ;
      RECT 0.8210 0.1330 0.8510 1.6120 ;
      RECT 3.1010 0.1330 3.1310 1.6120 ;
      RECT 2.9490 0.1340 2.9790 1.6120 ;
      RECT 2.7970 0.1330 2.8270 1.6120 ;
      RECT 2.6450 0.1330 2.6750 1.6120 ;
      RECT 3.2530 0.1330 3.2830 1.6120 ;
  END
END LSDNENSSX4_LVT

MACRO LSDNENSSX8_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.408 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0030 0.7650 4.1590 0.8150 ;
        RECT 4.0030 0.8150 4.0530 0.8890 ;
        RECT 4.0290 0.7050 4.1590 0.7650 ;
    END
    ANTENNAGATEAREA 0.0237 ;
  END EN

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.4080 0.0300 ;
        RECT 4.0790 0.0300 4.1290 0.4610 ;
        RECT 3.4710 0.0300 3.5210 0.3680 ;
        RECT 3.1670 0.0300 3.2170 0.3680 ;
        RECT 2.8630 0.0300 2.9130 0.3680 ;
        RECT 2.5590 0.0300 2.6090 0.3680 ;
    END
  END VSS

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.4080 1.7020 ;
        RECT 1.0390 1.3680 1.0890 1.6420 ;
        RECT 3.3190 1.0100 3.3690 1.6420 ;
        RECT 3.0150 1.1830 3.0650 1.6420 ;
        RECT 2.7110 1.1830 2.7610 1.6420 ;
        RECT 2.1030 1.3180 2.1530 1.6420 ;
        RECT 1.7990 1.3200 1.8490 1.6420 ;
        RECT 1.4950 1.3210 1.5450 1.6420 ;
        RECT 1.1910 1.3210 1.2410 1.6420 ;
        RECT 4.0780 1.0530 4.1280 1.6420 ;
        RECT 0.7350 1.3710 0.7850 1.6420 ;
        RECT 0.4310 1.3390 0.4810 1.6420 ;
        RECT 2.4070 1.3180 2.4570 1.6420 ;
    END
  END VDDL

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.8570 0.5110 0.9070 ;
        RECT 0.4010 0.9070 0.5110 0.9670 ;
    END
    ANTENNAGATEAREA 0.0237 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3430 0.8040 3.7510 0.8540 ;
        RECT 3.5880 0.8540 3.7510 0.9670 ;
        RECT 3.7010 0.5910 3.7510 0.8040 ;
        RECT 3.1670 0.8540 3.2170 1.5520 ;
        RECT 2.8630 0.8540 2.9130 1.5520 ;
        RECT 2.2550 0.8540 2.3050 1.0570 ;
        RECT 1.9510 0.8540 2.0010 1.0600 ;
        RECT 1.6470 0.8540 1.6970 1.0650 ;
        RECT 1.3430 0.8540 1.3930 1.0490 ;
        RECT 2.5590 0.8540 2.6090 1.5520 ;
        RECT 1.3430 0.5460 3.7510 0.5910 ;
        RECT 1.3430 0.5410 3.7450 0.5460 ;
        RECT 2.2550 0.1940 2.3050 0.5410 ;
        RECT 1.9510 0.1940 2.0010 0.5410 ;
        RECT 1.6470 0.1940 1.6970 0.5410 ;
        RECT 1.3430 0.1940 1.3930 0.5410 ;
    END
    ANTENNADIFFAREA 0.888 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 4.5230 1.7730 ;
    LAYER M1 ;
      RECT 3.8390 0.9810 3.9770 1.0310 ;
      RECT 3.9270 1.0310 3.9770 1.3200 ;
      RECT 3.8390 0.6500 3.9770 0.7000 ;
      RECT 3.5140 1.3200 3.9770 1.3700 ;
      RECT 3.9270 0.1950 3.9770 0.6500 ;
      RECT 3.9270 1.3700 3.9770 1.5200 ;
      RECT 3.8390 0.7000 3.8890 0.9810 ;
      RECT 1.0820 0.6610 2.3970 0.7110 ;
      RECT 1.0820 0.7110 1.1320 0.8040 ;
      RECT 1.0820 0.5820 1.1320 0.6610 ;
      RECT 0.8870 0.8040 1.1320 0.8540 ;
      RECT 0.8870 0.5320 1.1320 0.5820 ;
      RECT 0.8870 0.8540 0.9370 1.0140 ;
      RECT 0.8870 0.1940 0.9370 0.5320 ;
      RECT 2.4070 0.4240 3.6730 0.4740 ;
      RECT 3.6230 0.1940 3.6730 0.4240 ;
      RECT 2.4070 0.1380 2.4570 0.4240 ;
      RECT 0.4310 0.0880 2.4570 0.1380 ;
      RECT 2.7110 0.1940 2.7610 0.4240 ;
      RECT 3.0150 0.1940 3.0650 0.4240 ;
      RECT 3.3190 0.1940 3.3690 0.4240 ;
      RECT 1.0390 0.1380 1.0890 0.3680 ;
      RECT 1.1910 0.1380 1.2410 0.4600 ;
      RECT 0.4310 0.1380 0.4810 0.4610 ;
      RECT 0.7350 0.1380 0.7850 0.3680 ;
      RECT 1.4950 0.1380 1.5450 0.4600 ;
      RECT 1.7990 0.1380 1.8490 0.4600 ;
      RECT 2.1030 0.1380 2.1530 0.4600 ;
      RECT 0.5830 0.7730 0.8250 0.8230 ;
      RECT 0.5830 0.8230 0.6330 1.2420 ;
      RECT 0.7750 0.7000 0.8250 0.7730 ;
      RECT 0.7750 0.6500 1.0290 0.7000 ;
      RECT 0.7750 0.5510 0.8250 0.6500 ;
      RECT 0.5830 0.5010 0.8250 0.5510 ;
      RECT 0.5830 0.1940 0.6330 0.5010 ;
      RECT 2.4670 0.6610 3.6400 0.7110 ;
      RECT 0.2390 0.6600 0.7250 0.7100 ;
      RECT 0.2790 0.1950 0.3290 0.6600 ;
      RECT 0.2390 0.9660 0.3290 1.0160 ;
      RECT 0.2790 1.0160 0.3290 1.5240 ;
      RECT 0.2390 0.7100 0.2890 0.9660 ;
    LAYER PO ;
      RECT 1.1250 0.1330 1.1550 1.6120 ;
      RECT 0.8210 0.1330 0.8510 1.6120 ;
      RECT 0.6690 0.1330 0.6990 1.6120 ;
      RECT 3.5570 0.1340 3.5870 1.6120 ;
      RECT 3.4050 0.1330 3.4350 1.6120 ;
      RECT 3.2530 0.1340 3.2830 1.6120 ;
      RECT 3.1010 0.1330 3.1310 1.6120 ;
      RECT 2.9490 0.1330 2.9790 1.6120 ;
      RECT 2.6450 0.1330 2.6750 1.6120 ;
      RECT 2.7970 0.1340 2.8270 1.6120 ;
      RECT 2.3410 0.1330 2.3710 1.6120 ;
      RECT 2.4930 0.1340 2.5230 1.6120 ;
      RECT 2.1890 0.1330 2.2190 1.6120 ;
      RECT 2.0370 0.1330 2.0670 1.6120 ;
      RECT 1.8850 0.1330 1.9150 1.6120 ;
      RECT 1.5810 0.1330 1.6110 1.6120 ;
      RECT 1.7330 0.1340 1.7630 1.6120 ;
      RECT 1.2770 0.1330 1.3070 1.6120 ;
      RECT 3.8610 0.1330 3.8910 1.6120 ;
      RECT 3.7090 0.1340 3.7390 1.6120 ;
      RECT 1.4290 0.1340 1.4590 1.6120 ;
      RECT 0.3650 0.1330 0.3950 1.6120 ;
      RECT 0.5170 0.1330 0.5470 1.6120 ;
      RECT 0.9730 0.1330 1.0030 1.6120 ;
      RECT 0.0610 0.1330 0.0910 1.6040 ;
      RECT 0.2130 0.1330 0.2430 1.6120 ;
      RECT 4.1650 0.1340 4.1950 1.6120 ;
      RECT 4.0130 0.1330 4.0430 1.6120 ;
  END
END LSDNENSSX8_LVT

MACRO LSDNENX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.128 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9420 1.0020 1.1330 1.1360 ;
    END
    ANTENNAGATEAREA 0.0171 ;
  END EN

  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 3.0100 2.1280 3.0700 ;
        RECT 1.4660 3.0700 1.5760 3.1430 ;
        RECT 1.4660 2.9360 1.5760 3.0100 ;
        RECT 1.1910 2.5200 1.2410 3.0100 ;
        RECT 0.8870 2.5250 0.9370 3.0100 ;
    END
  END VDDH

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.1280 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.8070 ;
        RECT 1.0390 0.0300 1.0890 0.3480 ;
        RECT 1.7990 0.0300 1.8490 0.4850 ;
        RECT 0.7050 0.0300 0.7550 0.2960 ;
        RECT 0.7050 0.2960 0.7850 0.3570 ;
        RECT 0.7350 0.3570 0.7850 0.5050 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 2.1280 3.3740 ;
    END
  END VDDL

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.1280 1.7020 ;
        RECT 1.4660 1.7020 1.5760 1.7750 ;
        RECT 1.4660 1.5680 1.5760 1.6420 ;
        RECT 1.0390 1.4420 1.0890 1.6420 ;
        RECT 0.7350 1.3270 0.7850 1.6420 ;
        RECT 1.7990 1.3030 1.8490 1.6420 ;
        RECT 1.0390 1.7020 1.0890 2.1290 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5830 0.2300 0.6330 0.6940 ;
        RECT 0.5380 0.6940 0.6820 0.7780 ;
        RECT 0.4310 0.7780 0.6820 0.8280 ;
        RECT 0.4310 0.2300 0.4810 0.7780 ;
        RECT 0.4810 0.8280 0.5310 1.1980 ;
        RECT 0.4310 1.1980 0.5310 1.2620 ;
        RECT 0.4310 1.2620 0.4810 1.4520 ;
    END
    ANTENNADIFFAREA 0.1672 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7940 2.2130 1.1600 2.2630 ;
        RECT 0.9970 2.2630 1.1600 2.3650 ;
    END
    ANTENNAGATEAREA 0.0261 ;
  END A
  OBS
    LAYER NWELL ;
      RECT -0.1150 3.2240 2.2430 3.4590 ;
      RECT -0.1150 2.3510 0.1150 3.2240 ;
      RECT 2.0130 2.3510 2.2430 3.2240 ;
      RECT 0.5750 2.2340 1.4250 2.7640 ;
      RECT -0.1150 -0.1150 2.2430 0.9930 ;
    LAYER M1 ;
      RECT 0.5830 1.2920 0.6330 1.5390 ;
      RECT 0.2790 1.5390 0.6340 1.5890 ;
      RECT 0.2790 1.2920 0.3290 1.5390 ;
      RECT 0.8110 0.8380 0.9370 0.8880 ;
      RECT 0.8870 0.1880 0.9370 0.8380 ;
      RECT 0.8110 1.2190 0.9370 1.2690 ;
      RECT 0.8870 1.2690 0.9370 1.5830 ;
      RECT 0.8110 0.8880 0.8610 1.1560 ;
      RECT 0.6370 1.1560 0.8610 1.2060 ;
      RECT 0.8110 1.2060 0.8610 1.2190 ;
      RECT 0.6750 2.4230 1.0890 2.4730 ;
      RECT 1.0390 2.4730 1.0890 2.6900 ;
      RECT 0.6750 2.2630 0.7250 2.4230 ;
      RECT 0.1860 2.2130 0.7250 2.2630 ;
      RECT 0.6750 2.1280 0.7250 2.2130 ;
      RECT 0.6750 2.0780 0.9370 2.1280 ;
      RECT 0.8870 1.9760 0.9370 2.0780 ;
      RECT 0.7350 2.4730 0.7850 2.6900 ;
      RECT 0.1870 0.9240 0.4210 0.9740 ;
    LAYER PO ;
      RECT 1.7330 0.0690 1.7630 2.7800 ;
      RECT 0.3650 0.0890 0.3950 2.7800 ;
      RECT 1.1250 0.0870 1.1550 2.7780 ;
      RECT 1.8850 0.0690 1.9150 2.7800 ;
      RECT 0.9730 0.0890 1.0030 1.6690 ;
      RECT 1.5810 0.0690 1.6110 2.7800 ;
      RECT 1.2770 0.0750 1.3070 2.7800 ;
      RECT 1.4290 0.0750 1.4590 2.7800 ;
      RECT 2.0370 0.0740 2.0670 2.7800 ;
      RECT 0.9730 1.9210 1.0030 2.7820 ;
      RECT 0.8210 0.0780 0.8510 2.7800 ;
      RECT 0.0610 0.0890 0.0910 2.7800 ;
      RECT 0.6690 0.0890 0.6990 2.7810 ;
      RECT 0.5170 0.0890 0.5470 2.7800 ;
      RECT 0.2130 0.0890 0.2430 2.7800 ;
  END
END LSDNENX1_LVT

MACRO LSDNENX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.28 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9420 1.0020 1.1330 1.1360 ;
    END
    ANTENNAGATEAREA 0.0171 ;
  END EN

  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 3.0100 2.2800 3.0700 ;
        RECT 1.3140 3.0700 1.4240 3.1430 ;
        RECT 1.3140 2.9360 1.4240 3.0100 ;
        RECT 1.0390 2.5250 1.0890 3.0100 ;
        RECT 1.3430 2.5200 1.3930 2.9360 ;
    END
  END VDDH

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.2800 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.8070 ;
        RECT 1.6470 0.0300 1.6970 0.3450 ;
        RECT 1.0390 0.0300 1.0890 0.3480 ;
        RECT 1.3430 0.0300 1.3930 0.3450 ;
        RECT 1.9510 0.0300 2.0010 0.4850 ;
        RECT 0.7050 0.0300 0.7550 0.2960 ;
        RECT 0.7050 0.2960 0.7850 0.3570 ;
        RECT 0.7350 0.3570 0.7850 0.5050 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 2.2800 3.3740 ;
    END
  END VDDL

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.2800 1.7020 ;
        RECT 1.9220 1.7020 2.0320 1.7750 ;
        RECT 1.9220 1.5680 2.0320 1.6420 ;
        RECT 1.0390 1.4420 1.0890 1.6420 ;
        RECT 1.6470 1.3630 1.6970 1.6420 ;
        RECT 1.3430 1.4420 1.3930 1.6420 ;
        RECT 0.7350 1.3270 0.7850 1.6420 ;
        RECT 1.0390 1.7020 1.0890 2.1290 ;
        RECT 1.9510 1.3480 2.0010 1.5680 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8660 0.6700 1.9160 0.6940 ;
        RECT 1.8660 0.6940 2.0590 0.8280 ;
        RECT 1.4950 0.6200 1.9160 0.6700 ;
        RECT 1.8660 0.8280 1.9160 1.1810 ;
        RECT 1.7990 0.2170 1.8490 0.6200 ;
        RECT 1.4950 0.1850 1.5450 0.6200 ;
        RECT 1.4950 1.1810 1.9160 1.2310 ;
        RECT 1.7990 1.2310 1.8490 1.5830 ;
        RECT 1.4950 1.2310 1.5450 1.5830 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9460 2.2130 1.3120 2.2630 ;
        RECT 1.1490 2.2630 1.3120 2.3650 ;
    END
    ANTENNAGATEAREA 0.0261 ;
  END A
  OBS
    LAYER NWELL ;
      RECT -0.1150 3.2240 2.3950 3.4590 ;
      RECT -0.1150 2.3510 0.1150 3.2240 ;
      RECT 2.1650 2.3510 2.3950 3.2240 ;
      RECT 0.5750 2.2340 1.6170 2.7640 ;
      RECT -0.1150 -0.1150 2.3950 0.9930 ;
    LAYER M1 ;
      RECT 1.2200 1.0280 1.3330 1.0780 ;
      RECT 0.5830 0.2300 0.6330 0.7720 ;
      RECT 0.4310 0.2300 0.4810 0.7720 ;
      RECT 0.4810 0.8220 0.5310 1.1980 ;
      RECT 0.4310 1.1980 0.5310 1.2620 ;
      RECT 0.4310 1.2620 0.4810 1.4520 ;
      RECT 1.2200 0.9510 1.2700 1.0280 ;
      RECT 1.0620 0.9010 1.2700 0.9510 ;
      RECT 1.0620 0.8220 1.1120 0.9010 ;
      RECT 0.4310 0.7720 1.1120 0.8220 ;
      RECT 1.3830 1.0330 1.7890 1.0830 ;
      RECT 1.1910 1.2510 1.2410 1.5830 ;
      RECT 1.3830 1.0830 1.4330 1.2010 ;
      RECT 1.3830 0.7050 1.4330 1.0330 ;
      RECT 1.1910 1.2010 1.4330 1.2510 ;
      RECT 1.1720 0.6550 1.4330 0.7050 ;
      RECT 0.8270 2.4230 1.2410 2.4730 ;
      RECT 1.1910 2.4730 1.2410 2.6900 ;
      RECT 0.8270 2.2850 0.8770 2.4230 ;
      RECT 0.7660 2.2630 0.8770 2.2850 ;
      RECT 0.1860 2.2130 0.8770 2.2630 ;
      RECT 0.7660 2.1840 0.8770 2.2130 ;
      RECT 0.8270 2.1280 0.8770 2.1840 ;
      RECT 0.8870 2.4730 0.9370 2.6900 ;
      RECT 0.8270 2.0780 0.9370 2.1280 ;
      RECT 0.8870 1.9760 0.9370 2.0780 ;
      RECT 0.2790 1.5340 0.6330 1.5840 ;
      RECT 0.5830 1.2920 0.6330 1.5340 ;
      RECT 0.2790 1.2920 0.3290 1.5340 ;
      RECT 0.8110 0.1880 0.9370 0.2380 ;
      RECT 0.8110 0.0880 0.8610 0.1880 ;
      RECT 0.8870 0.2380 0.9370 0.4210 ;
      RECT 0.8110 1.2190 0.9370 1.2690 ;
      RECT 0.8870 1.2690 0.9370 1.5830 ;
      RECT 0.6370 1.1560 0.8610 1.2060 ;
      RECT 0.8110 1.2060 0.8610 1.2190 ;
      RECT 0.8110 1.1400 0.8610 1.1560 ;
      RECT 0.1870 0.9240 0.4210 0.9740 ;
    LAYER PO ;
      RECT 1.8850 0.0690 1.9150 2.7800 ;
      RECT 0.3650 0.0890 0.3950 2.7800 ;
      RECT 1.1250 0.0870 1.1550 2.7780 ;
      RECT 2.0370 0.0690 2.0670 2.7800 ;
      RECT 0.9730 0.0890 1.0030 1.6690 ;
      RECT 1.5810 0.0660 1.6110 2.7800 ;
      RECT 1.2770 0.0750 1.3070 2.7800 ;
      RECT 1.4290 0.0750 1.4590 2.7800 ;
      RECT 2.1890 0.0740 2.2190 2.7800 ;
      RECT 1.7330 0.0660 1.7630 2.7800 ;
      RECT 0.9730 1.9210 1.0030 2.7820 ;
      RECT 0.8210 0.0880 0.8510 2.7800 ;
      RECT 0.0610 0.0890 0.0910 2.7800 ;
      RECT 0.6690 0.0890 0.6990 2.7810 ;
      RECT 0.5170 0.0890 0.5470 2.7800 ;
      RECT 0.2130 0.0890 0.2430 2.7800 ;
  END
END LSDNENX2_LVT

MACRO LSDNENX4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.584 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9420 1.0020 1.1330 1.1360 ;
    END
    ANTENNAGATEAREA 0.0171 ;
  END EN

  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 3.0100 2.5840 3.0700 ;
        RECT 1.3140 3.0700 1.4240 3.1430 ;
        RECT 1.3140 2.9360 1.4240 3.0100 ;
        RECT 1.0390 2.5250 1.0890 3.0100 ;
        RECT 1.3430 2.5200 1.3930 2.9360 ;
    END
  END VDDH

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.5840 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.8070 ;
        RECT 1.6470 0.0300 1.6970 0.3450 ;
        RECT 1.0390 0.0300 1.0890 0.3480 ;
        RECT 1.9510 0.0300 2.0010 0.3450 ;
        RECT 1.3430 0.0300 1.3930 0.3450 ;
        RECT 2.2550 0.0300 2.3050 0.4850 ;
        RECT 0.7050 0.0300 0.7550 0.3430 ;
        RECT 0.7050 0.3430 0.7850 0.4040 ;
        RECT 0.7350 0.4040 0.7850 0.5870 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 2.5840 3.3740 ;
    END
  END VDDL

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.5840 1.7020 ;
        RECT 2.2260 1.7020 2.3360 1.7750 ;
        RECT 2.2260 1.5680 2.3360 1.6420 ;
        RECT 1.0390 1.4420 1.0890 1.6420 ;
        RECT 1.6470 1.3630 1.6970 1.6420 ;
        RECT 1.9510 1.3630 2.0010 1.6420 ;
        RECT 1.3430 1.4420 1.3930 1.6420 ;
        RECT 0.7350 1.3270 0.7850 1.6420 ;
        RECT 1.0390 1.7020 1.0890 2.1290 ;
        RECT 2.2550 1.3170 2.3050 1.5680 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2120 0.6700 2.2620 0.6940 ;
        RECT 2.2120 0.6940 2.3630 0.8280 ;
        RECT 1.4950 0.6200 2.2620 0.6700 ;
        RECT 2.2120 0.8280 2.2620 1.2010 ;
        RECT 2.1030 0.2170 2.1530 0.6200 ;
        RECT 1.7990 0.2170 1.8490 0.6200 ;
        RECT 1.4950 0.1850 1.5450 0.6200 ;
        RECT 1.4950 1.2010 2.2620 1.2510 ;
        RECT 2.1030 1.2510 2.1530 1.5830 ;
        RECT 1.4950 1.2510 1.5450 1.5830 ;
        RECT 1.7990 1.2510 1.8490 1.5830 ;
    END
    ANTENNADIFFAREA 0.3976 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9460 2.2130 1.3120 2.2630 ;
        RECT 1.1490 2.2630 1.3120 2.3650 ;
    END
    ANTENNAGATEAREA 0.0261 ;
  END A
  OBS
    LAYER NWELL ;
      RECT -0.1150 3.2240 2.6990 3.4590 ;
      RECT -0.1150 2.3510 0.1150 3.2240 ;
      RECT 2.4690 2.3510 2.6990 3.2240 ;
      RECT 0.5750 2.2340 1.6170 2.7640 ;
      RECT -0.1150 -0.1150 2.6990 0.9930 ;
    LAYER M1 ;
      RECT 1.2200 1.0280 1.3330 1.0780 ;
      RECT 0.5830 0.2300 0.6330 0.7720 ;
      RECT 0.4310 0.2300 0.4810 0.7720 ;
      RECT 0.4810 0.8220 0.5310 1.1980 ;
      RECT 0.4310 1.1980 0.5310 1.2620 ;
      RECT 0.4310 1.2620 0.4810 1.4520 ;
      RECT 1.2200 0.9510 1.2700 1.0280 ;
      RECT 1.0620 0.9010 1.2700 0.9510 ;
      RECT 1.0620 0.8220 1.1120 0.9010 ;
      RECT 0.4310 0.7720 1.1120 0.8220 ;
      RECT 1.3830 1.0330 2.1240 1.0830 ;
      RECT 1.1910 1.2510 1.2410 1.5830 ;
      RECT 1.3830 1.0830 1.4330 1.2010 ;
      RECT 1.3830 0.8510 1.4330 1.0330 ;
      RECT 1.1910 1.2010 1.4330 1.2510 ;
      RECT 1.1720 0.8010 1.4330 0.8510 ;
      RECT 0.8270 2.4230 1.2410 2.4730 ;
      RECT 1.1910 2.4730 1.2410 2.6900 ;
      RECT 0.8270 2.2850 0.8770 2.4230 ;
      RECT 0.7660 2.2630 0.8770 2.2850 ;
      RECT 0.1860 2.2130 0.8770 2.2630 ;
      RECT 0.7660 2.1840 0.8770 2.2130 ;
      RECT 0.8270 2.1280 0.8770 2.1840 ;
      RECT 0.8870 2.4730 0.9370 2.6900 ;
      RECT 0.8270 2.0780 0.9370 2.1280 ;
      RECT 0.8870 1.9760 0.9370 2.0780 ;
      RECT 0.2790 1.5340 0.6330 1.5840 ;
      RECT 0.5830 1.2920 0.6330 1.5340 ;
      RECT 0.2790 1.2920 0.3290 1.5340 ;
      RECT 0.8110 0.1880 0.9370 0.2380 ;
      RECT 0.8110 0.0880 0.8610 0.1880 ;
      RECT 0.8870 0.2380 0.9370 0.4210 ;
      RECT 0.8110 1.2190 0.9370 1.2690 ;
      RECT 0.8870 1.2690 0.9370 1.5830 ;
      RECT 0.6370 1.1560 0.8610 1.2060 ;
      RECT 0.8110 1.2060 0.8610 1.2190 ;
      RECT 0.8110 1.1400 0.8610 1.1560 ;
      RECT 0.1870 0.9240 0.4210 0.9740 ;
    LAYER PO ;
      RECT 2.0370 0.0620 2.0670 2.7800 ;
      RECT 2.1890 0.0620 2.2190 2.7800 ;
      RECT 0.3650 0.0890 0.3950 2.7800 ;
      RECT 1.1250 0.0870 1.1550 2.7780 ;
      RECT 2.3410 0.0620 2.3710 2.7800 ;
      RECT 1.8850 0.0620 1.9150 2.7800 ;
      RECT 0.9730 0.0890 1.0030 1.6690 ;
      RECT 1.5810 0.0620 1.6110 2.7800 ;
      RECT 1.2770 0.0680 1.3070 2.7800 ;
      RECT 1.4290 0.0680 1.4590 2.7800 ;
      RECT 2.4930 0.0670 2.5230 2.7800 ;
      RECT 1.7330 0.0620 1.7630 2.7800 ;
      RECT 0.9730 1.9210 1.0030 2.7820 ;
      RECT 0.8210 0.0780 0.8510 2.7800 ;
      RECT 0.0610 0.0890 0.0910 2.7800 ;
      RECT 0.6690 0.0890 0.6990 2.7810 ;
      RECT 0.5170 0.0890 0.5470 2.7800 ;
      RECT 0.2130 0.0890 0.2430 2.7800 ;
  END
END LSDNENX4_LVT

MACRO LSDNENX8_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.344 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9420 1.0020 1.1330 1.1360 ;
    END
    ANTENNAGATEAREA 0.0171 ;
  END EN

  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 3.0100 3.3440 3.0700 ;
        RECT 1.9220 3.0700 2.0320 3.1430 ;
        RECT 1.9220 2.9360 2.0320 3.0100 ;
        RECT 1.3430 2.5200 1.3930 3.0100 ;
        RECT 1.0390 2.5250 1.0890 3.0100 ;
    END
  END VDDH

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.3440 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.8070 ;
        RECT 2.7110 0.0300 2.7610 0.3450 ;
        RECT 1.7990 0.0300 1.8490 0.3450 ;
        RECT 1.0390 0.0300 1.0890 0.3480 ;
        RECT 2.4070 0.0300 2.4570 0.3500 ;
        RECT 2.1030 0.0300 2.1530 0.3450 ;
        RECT 1.1910 0.0300 1.2410 0.3450 ;
        RECT 1.4950 0.0300 1.5450 0.3450 ;
        RECT 3.0150 0.0300 3.0650 0.4850 ;
        RECT 0.7050 0.0300 0.7550 0.3430 ;
        RECT 0.7050 0.3430 0.7850 0.4040 ;
        RECT 0.7350 0.4040 0.7850 0.5870 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 3.3440 3.3740 ;
    END
  END VDDL

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.3440 1.7020 ;
        RECT 2.9860 1.7020 3.0960 1.7750 ;
        RECT 2.9860 1.5680 3.0960 1.6420 ;
        RECT 1.0390 1.7020 1.0890 2.1290 ;
        RECT 1.0390 1.4420 1.0890 1.6420 ;
        RECT 2.7110 1.3630 2.7610 1.6420 ;
        RECT 1.7990 1.3630 1.8490 1.6420 ;
        RECT 2.4070 1.3630 2.4570 1.6420 ;
        RECT 2.1030 1.3630 2.1530 1.6420 ;
        RECT 1.1910 1.4420 1.2410 1.6420 ;
        RECT 1.4950 1.4420 1.5450 1.6420 ;
        RECT 0.7350 1.3270 0.7850 1.6420 ;
        RECT 3.0150 1.3380 3.0650 1.5680 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9300 0.6700 2.9800 0.6940 ;
        RECT 2.9300 0.6940 3.1230 0.8280 ;
        RECT 1.6470 0.6200 2.9800 0.6700 ;
        RECT 2.9300 0.8280 2.9800 1.1750 ;
        RECT 2.8630 0.2170 2.9130 0.6200 ;
        RECT 2.2550 0.2170 2.3050 0.6200 ;
        RECT 2.5590 0.1850 2.6090 0.6200 ;
        RECT 1.9510 0.2170 2.0010 0.6200 ;
        RECT 1.6470 0.1850 1.6970 0.6200 ;
        RECT 1.6470 1.1750 2.9800 1.2250 ;
        RECT 2.5590 1.2250 2.6090 1.4150 ;
        RECT 2.8630 1.2250 2.9130 1.4150 ;
        RECT 2.2550 1.2250 2.3050 1.4140 ;
        RECT 1.6470 1.2250 1.6970 1.4130 ;
        RECT 1.9510 1.2250 2.0010 1.4130 ;
    END
    ANTENNADIFFAREA 0.6952 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9460 2.2130 1.3120 2.2630 ;
        RECT 1.1490 2.2630 1.3120 2.3650 ;
    END
    ANTENNAGATEAREA 0.0261 ;
  END A
  OBS
    LAYER NWELL ;
      RECT -0.1150 3.2240 3.4590 3.4590 ;
      RECT -0.1150 2.3510 0.1150 3.2240 ;
      RECT 3.2290 2.3510 3.4590 3.2240 ;
      RECT 0.5750 2.2340 1.6170 2.7640 ;
      RECT -0.1150 -0.1150 3.4590 0.9930 ;
    LAYER M1 ;
      RECT 1.5350 1.0330 2.8630 1.0830 ;
      RECT 1.5350 0.8510 1.5850 1.0330 ;
      RECT 1.5350 1.0830 1.5850 1.2010 ;
      RECT 1.3430 0.8010 1.5850 0.8510 ;
      RECT 1.3430 1.2010 1.5850 1.2510 ;
      RECT 1.3430 0.8510 1.3930 0.9170 ;
      RECT 1.3430 1.2510 1.3930 1.3250 ;
      RECT 1.2200 1.0280 1.4850 1.0780 ;
      RECT 0.5830 0.2300 0.6330 0.7720 ;
      RECT 0.4310 0.2300 0.4810 0.7720 ;
      RECT 0.4810 0.8220 0.5310 1.1980 ;
      RECT 0.4310 1.1980 0.5310 1.2620 ;
      RECT 0.4310 1.2620 0.4810 1.4520 ;
      RECT 1.2200 0.8220 1.2700 1.0280 ;
      RECT 0.4310 0.7720 1.2700 0.8220 ;
      RECT 0.8270 2.4230 1.2410 2.4730 ;
      RECT 1.1910 2.4730 1.2410 2.6900 ;
      RECT 0.8270 2.2850 0.8770 2.4230 ;
      RECT 0.7660 2.2630 0.8770 2.2850 ;
      RECT 0.1860 2.2130 0.8770 2.2630 ;
      RECT 0.7660 2.1840 0.8770 2.2130 ;
      RECT 0.8270 2.1280 0.8770 2.1840 ;
      RECT 0.8870 2.4730 0.9370 2.6900 ;
      RECT 0.8270 2.0780 0.9370 2.1280 ;
      RECT 0.8870 1.9760 0.9370 2.0780 ;
      RECT 0.1870 0.9240 0.4210 0.9740 ;
      RECT 0.2790 1.5340 0.6330 1.5840 ;
      RECT 0.5830 1.2920 0.6330 1.5340 ;
      RECT 0.2790 1.2920 0.3290 1.5340 ;
      RECT 0.8110 0.1880 0.9370 0.2380 ;
      RECT 0.8110 0.0880 0.8610 0.1880 ;
      RECT 0.8870 0.2380 0.9370 0.4210 ;
      RECT 0.8110 1.2190 0.9370 1.2690 ;
      RECT 0.8870 1.2690 0.9370 1.5830 ;
      RECT 0.6370 1.1560 0.8610 1.2060 ;
      RECT 0.8110 1.2060 0.8610 1.2190 ;
      RECT 0.8110 1.1400 0.8610 1.1560 ;
    LAYER PO ;
      RECT 3.2530 0.0730 3.2830 2.7800 ;
      RECT 2.0370 0.0680 2.0670 2.7800 ;
      RECT 2.1890 0.0680 2.2190 2.7800 ;
      RECT 2.3410 0.0680 2.3710 2.7800 ;
      RECT 2.4930 0.0680 2.5230 2.7800 ;
      RECT 2.6450 0.0680 2.6750 2.7800 ;
      RECT 2.7970 0.0680 2.8270 2.7800 ;
      RECT 0.3650 0.0890 0.3950 2.7800 ;
      RECT 1.1250 0.0870 1.1550 2.7780 ;
      RECT 2.9490 0.0680 2.9790 2.7800 ;
      RECT 1.8850 0.0680 1.9150 2.7800 ;
      RECT 0.9730 0.0890 1.0030 1.6690 ;
      RECT 1.5810 0.0680 1.6110 2.7800 ;
      RECT 1.2770 0.0680 1.3070 2.7800 ;
      RECT 1.4290 0.0680 1.4590 2.7800 ;
      RECT 3.1010 0.0730 3.1310 2.7800 ;
      RECT 1.7330 0.0680 1.7630 2.7800 ;
      RECT 0.9730 1.9210 1.0030 2.7820 ;
      RECT 0.8210 0.0880 0.8510 2.7800 ;
      RECT 0.0610 0.0890 0.0910 2.7800 ;
      RECT 0.6690 0.0890 0.6990 2.7810 ;
      RECT 0.5170 0.0890 0.5470 2.7800 ;
      RECT 0.2130 0.0890 0.2430 2.7800 ;
  END
END LSDNENX8_LVT

MACRO LSDNSSX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.064 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6750 0.4210 0.7250 ;
        RECT 0.2490 0.7250 0.3620 0.8150 ;
    END
    ANTENNAGATEAREA 0.012 ;
  END A

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.0640 1.7020 ;
        RECT 0.2790 0.8750 0.3290 1.6420 ;
        RECT 0.7350 0.9120 0.7850 1.6420 ;
    END
  END VDDL

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.0640 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.5480 ;
        RECT 0.7350 0.0300 0.7850 0.4870 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5830 0.8120 0.8410 0.8620 ;
        RECT 0.5830 0.8620 0.6330 1.5460 ;
        RECT 0.7910 0.6630 0.8410 0.8120 ;
        RECT 0.7910 0.5870 0.9670 0.6630 ;
        RECT 0.5830 0.5370 0.9670 0.5870 ;
        RECT 0.5830 0.3350 0.6330 0.5370 ;
    END
    ANTENNADIFFAREA 0.1081 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.1790 1.7730 ;
    LAYER M1 ;
      RECT 0.4910 0.6600 0.7250 0.7100 ;
      RECT 0.4560 0.8870 0.5210 0.9370 ;
      RECT 0.4310 0.8870 0.4810 1.0610 ;
      RECT 0.4310 0.8870 0.4740 0.9370 ;
      RECT 0.4310 0.4660 0.4810 0.5710 ;
      RECT 0.4710 0.4660 0.5210 0.9370 ;
    LAYER PO ;
      RECT 0.0610 0.0710 0.0910 1.6060 ;
      RECT 0.3650 0.0690 0.3950 1.6060 ;
      RECT 0.2130 0.0710 0.2430 1.6060 ;
      RECT 0.5170 0.0710 0.5470 1.6060 ;
      RECT 0.6690 0.0690 0.6990 1.6060 ;
      RECT 0.9730 0.0710 1.0030 1.6060 ;
      RECT 0.8210 0.0710 0.8510 1.6060 ;
  END
END LSDNSSX1_LVT

MACRO LSDNSSX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.216 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6750 0.4210 0.7250 ;
        RECT 0.2490 0.7250 0.3620 0.8150 ;
    END
    ANTENNAGATEAREA 0.0255 ;
  END A

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.2160 1.7020 ;
        RECT 0.2790 0.8730 0.3290 1.6420 ;
        RECT 0.7350 0.9120 0.7850 1.6420 ;
    END
  END VDDL

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.2160 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.5480 ;
        RECT 0.7350 0.0300 0.7850 0.4870 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5830 0.8120 0.9930 0.8620 ;
        RECT 0.5830 0.8620 0.6330 1.5460 ;
        RECT 0.8870 0.8620 0.9370 1.5460 ;
        RECT 0.9430 0.6630 0.9930 0.8120 ;
        RECT 0.9430 0.5870 1.1190 0.6630 ;
        RECT 0.5830 0.5370 1.1190 0.5870 ;
        RECT 0.5830 0.3350 0.6330 0.5370 ;
        RECT 0.8870 0.3350 0.9370 0.5370 ;
    END
    ANTENNADIFFAREA 0.2162 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.3310 1.7730 ;
    LAYER M1 ;
      RECT 0.4910 0.6600 0.8770 0.7100 ;
      RECT 0.4560 0.8870 0.5210 0.9370 ;
      RECT 0.4310 0.8870 0.4810 1.3370 ;
      RECT 0.4310 0.3740 0.4810 0.5480 ;
      RECT 0.4710 0.4660 0.5210 0.9370 ;
    LAYER PO ;
      RECT 0.0610 0.0710 0.0910 1.6060 ;
      RECT 0.3650 0.0690 0.3950 1.6060 ;
      RECT 0.2130 0.0710 0.2430 1.6060 ;
      RECT 1.1250 0.0710 1.1550 1.6060 ;
      RECT 0.5170 0.0710 0.5470 1.6060 ;
      RECT 0.6690 0.0690 0.6990 1.6060 ;
      RECT 0.9730 0.0710 1.0030 1.6060 ;
      RECT 0.8210 0.0710 0.8510 1.6060 ;
  END
END LSDNSSX2_LVT

MACRO LSDNSSX4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.52 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6600 0.4210 0.7100 ;
        RECT 0.2490 0.7100 0.3620 0.8150 ;
    END
    ANTENNAGATEAREA 0.0318 ;
  END A

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.5200 1.7020 ;
        RECT 1.0390 0.9120 1.0890 1.6420 ;
        RECT 0.2790 0.8690 0.3290 1.6420 ;
        RECT 0.7350 0.9120 0.7850 1.6420 ;
    END
  END VDDL

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.5200 0.0300 ;
        RECT 1.0390 0.0300 1.0890 0.4870 ;
        RECT 0.2790 0.0300 0.3290 0.5510 ;
        RECT 0.7350 0.0300 0.7850 0.4870 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5830 0.8120 1.2970 0.8620 ;
        RECT 1.1910 0.8620 1.2410 1.5460 ;
        RECT 0.5830 0.8620 0.6330 1.5460 ;
        RECT 0.8870 0.8620 0.9370 1.5460 ;
        RECT 1.2470 0.6630 1.2970 0.8120 ;
        RECT 1.2470 0.5870 1.4230 0.6630 ;
        RECT 0.5830 0.5370 1.4230 0.5870 ;
        RECT 0.5830 0.3350 0.6330 0.5370 ;
        RECT 1.1910 0.3350 1.2410 0.5370 ;
        RECT 0.8870 0.3350 0.9370 0.5370 ;
    END
    ANTENNADIFFAREA 0.3456 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.6350 1.7730 ;
    LAYER M1 ;
      RECT 0.4910 0.6600 1.1810 0.7100 ;
      RECT 0.4560 0.8870 0.5210 0.9370 ;
      RECT 0.4310 0.8870 0.4810 1.5210 ;
      RECT 0.4310 0.3770 0.4810 0.5510 ;
      RECT 0.4710 0.4660 0.5210 0.9370 ;
    LAYER PO ;
      RECT 0.0610 0.0710 0.0910 1.6060 ;
      RECT 0.3650 0.0690 0.3950 1.6060 ;
      RECT 0.2130 0.0710 0.2430 1.6060 ;
      RECT 1.1250 0.0710 1.1550 1.6060 ;
      RECT 0.5170 0.0710 0.5470 1.6060 ;
      RECT 0.6690 0.0690 0.6990 1.6060 ;
      RECT 0.9730 0.0710 1.0030 1.6060 ;
      RECT 0.8210 0.0710 0.8510 1.6060 ;
      RECT 1.2770 0.0710 1.3070 1.6060 ;
      RECT 1.4290 0.0710 1.4590 1.6060 ;
  END
END LSDNSSX4_LVT

MACRO LASRX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9470 0.7880 1.1190 0.9670 ;
    END
    ANTENNAGATEAREA 0.0261 ;
  END D

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.8000 0.0300 ;
        RECT 2.8630 0.0300 2.9130 0.2200 ;
        RECT 0.4310 0.0300 0.4810 0.4500 ;
        RECT 0.5830 0.0300 0.6330 0.4500 ;
        RECT 3.4710 0.0300 3.5210 0.2200 ;
        RECT 3.1670 0.0300 3.2170 0.2200 ;
        RECT 2.7110 0.0300 2.7610 0.2440 ;
        RECT 0.8870 0.2440 2.7610 0.2940 ;
        RECT 0.8870 0.2940 0.9370 0.4210 ;
        RECT 2.7110 0.2940 2.7610 0.3540 ;
    END
  END VSS

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0150 0.1480 3.0650 0.3950 ;
        RECT 3.0150 0.3950 3.5610 0.4450 ;
        RECT 3.5110 0.4450 3.5610 1.0090 ;
        RECT 3.0150 1.0090 3.5610 1.0590 ;
        RECT 3.2890 1.0590 3.3990 1.1190 ;
        RECT 3.0150 1.0590 3.0650 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.8000 1.7020 ;
        RECT 2.8630 1.1700 2.9130 1.6420 ;
        RECT 3.4710 1.3570 3.5210 1.6420 ;
        RECT 3.1670 1.1700 3.2170 1.6420 ;
        RECT 0.4910 1.3540 0.5410 1.6420 ;
        RECT 2.7510 1.3780 2.8010 1.6420 ;
        RECT 0.4310 1.3040 1.1050 1.3540 ;
        RECT 2.1280 1.3280 2.8010 1.3780 ;
        RECT 0.4310 1.0880 0.4810 1.3040 ;
        RECT 0.5830 1.1010 0.6330 1.3040 ;
        RECT 2.1280 1.2430 2.1780 1.3280 ;
        RECT 1.7830 1.1930 2.1780 1.2430 ;
    END
  END VDD

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7690 1.3130 1.9230 1.4230 ;
    END
    ANTENNAGATEAREA 0.0261 ;
  END SETB

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.3030 0.2950 3.6610 0.3450 ;
        RECT 3.6110 0.3450 3.6610 1.2210 ;
        RECT 3.3190 1.2210 3.6610 1.2710 ;
        RECT 3.4460 1.1610 3.5560 1.2210 ;
        RECT 3.3190 1.2710 3.3690 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 1.4240 0.4210 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0990 0.5530 1.2710 0.6660 ;
    END
    ANTENNAGATEAREA 0.0441 ;
  END RSTB
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 3.9150 1.7730 ;
      RECT 0.5320 0.6660 0.8360 0.6790 ;
    LAYER M1 ;
      RECT 1.9510 0.6040 3.1570 0.6540 ;
      RECT 1.9510 0.4800 2.0010 0.6040 ;
      RECT 2.2950 0.6540 2.3450 0.8780 ;
      RECT 1.6300 0.8780 2.3450 0.9280 ;
      RECT 1.4550 0.6060 1.5450 0.6560 ;
      RECT 1.4950 0.4300 1.5450 0.6060 ;
      RECT 1.4550 0.6560 1.5050 1.0010 ;
      RECT 1.4950 0.3800 2.1530 0.4300 ;
      RECT 1.4550 1.0010 2.1740 1.0510 ;
      RECT 2.1030 0.4300 2.1530 0.5540 ;
      RECT 1.7980 0.4300 1.8480 0.6180 ;
      RECT 1.7070 0.6180 1.8480 0.6680 ;
      RECT 2.0100 1.4280 2.2450 1.4780 ;
      RECT 1.1750 0.4180 1.3930 0.4680 ;
      RECT 1.3430 0.4680 1.3930 1.3080 ;
      RECT 1.1910 1.3080 1.3930 1.3580 ;
      RECT 1.1910 1.2160 1.2410 1.3080 ;
      RECT 0.8700 1.1660 1.2410 1.2160 ;
      RECT 0.7350 0.0960 2.1240 0.1460 ;
      RECT 0.7350 0.5180 0.8610 0.5680 ;
      RECT 0.8110 0.5680 0.8610 0.7180 ;
      RECT 0.7350 0.7180 0.8610 0.7680 ;
      RECT 0.7350 0.1460 0.7850 0.5180 ;
      RECT 0.7350 0.7680 0.7850 0.9140 ;
      RECT 0.2790 0.6180 0.7250 0.6680 ;
      RECT 0.2790 0.6680 0.3290 1.3540 ;
      RECT 0.2790 0.4220 0.3290 0.6180 ;
      RECT 3.2430 0.6040 3.4610 0.6540 ;
      RECT 3.2430 0.5450 3.2930 0.6040 ;
      RECT 3.2430 0.6540 3.2930 0.8060 ;
      RECT 2.2390 0.4950 3.2930 0.5450 ;
      RECT 2.7270 0.8060 3.2930 0.8560 ;
      RECT 2.7270 0.8560 2.7770 1.1180 ;
      RECT 2.2390 1.1180 2.7770 1.1680 ;
      RECT 1.5550 0.7180 2.2450 0.7680 ;
      RECT 1.0990 1.5280 2.7010 1.5780 ;
      RECT 0.6590 1.4280 1.6370 1.4780 ;
      RECT 0.6590 1.4780 0.7090 1.5840 ;
    LAYER PO ;
      RECT 3.7090 0.0680 3.7390 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 1.2770 0.0680 1.3070 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 2.1890 0.9320 2.2190 1.6060 ;
      RECT 1.4290 0.0680 1.4590 0.6420 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 2.1890 0.0680 2.2190 0.7960 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 1.4290 0.8820 1.4590 1.6060 ;
  END
END LASRX2_LVT

MACRO LASX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.192 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9470 0.6660 1.1190 0.8150 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END D

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.1920 0.0300 ;
        RECT 2.7110 0.0300 2.7610 0.2200 ;
        RECT 0.5830 0.0300 0.6330 0.4500 ;
        RECT 0.4310 0.0300 0.4810 0.4500 ;
        RECT 2.4070 0.0300 2.4570 0.2880 ;
        RECT 0.8870 0.2880 2.4570 0.3380 ;
        RECT 0.8870 0.3380 0.9370 0.4620 ;
    END
  END VSS

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5590 1.0690 2.9430 1.1190 ;
        RECT 2.8330 1.0090 2.9430 1.0690 ;
        RECT 2.5590 1.1190 2.6090 1.5460 ;
        RECT 2.8930 0.3590 2.9430 1.0090 ;
        RECT 2.5590 0.3090 2.9430 0.3590 ;
        RECT 2.5590 0.1480 2.6090 0.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.1920 1.7020 ;
        RECT 2.7110 1.1700 2.7610 1.6420 ;
        RECT 0.5590 1.1270 0.6090 1.6420 ;
        RECT 2.4230 1.3780 2.4730 1.6420 ;
        RECT 0.4310 1.0770 0.9370 1.1270 ;
        RECT 1.9760 1.3280 2.4730 1.3780 ;
        RECT 0.4310 0.8610 0.4810 1.0770 ;
        RECT 0.5830 0.8740 0.6330 1.0770 ;
        RECT 0.8870 1.1270 0.9370 1.3430 ;
        RECT 1.9760 1.3150 2.0260 1.3280 ;
        RECT 1.6310 1.2650 2.0260 1.3150 ;
    END
  END VDD

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6170 1.4650 1.7710 1.5750 ;
    END
    ANTENNAGATEAREA 0.018 ;
  END SETB

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9850 1.1610 3.0960 1.2210 ;
        RECT 2.8630 1.2210 3.0960 1.2710 ;
        RECT 3.0450 0.2040 3.0950 1.1610 ;
        RECT 2.8630 1.2710 2.9130 1.5460 ;
        RECT 2.8470 0.1540 3.0950 0.2040 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 1.3130 0.4050 1.4230 ;
        RECT 0.3550 1.4230 0.4050 1.5840 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 3.3070 1.7730 ;
      RECT 0.2180 0.6680 0.8410 0.6790 ;
    LAYER M1 ;
      RECT 1.7990 0.6040 2.7010 0.6540 ;
      RECT 1.7990 0.5100 1.8490 0.6040 ;
      RECT 2.1430 0.6540 2.1930 1.0650 ;
      RECT 1.4790 1.0650 2.1930 1.1150 ;
      RECT 1.5550 0.6180 1.6960 0.6680 ;
      RECT 1.6460 0.4600 1.6960 0.6180 ;
      RECT 1.3430 0.4100 2.0170 0.4600 ;
      RECT 1.3430 0.4600 1.3930 0.6060 ;
      RECT 1.3030 0.6060 1.3930 0.6560 ;
      RECT 1.3030 0.6560 1.3530 1.1650 ;
      RECT 1.3030 1.1650 2.0220 1.2150 ;
      RECT 0.7350 0.0960 1.9720 0.1460 ;
      RECT 0.7350 0.5180 0.8610 0.5680 ;
      RECT 0.8110 0.5680 0.8610 0.7180 ;
      RECT 0.7350 0.7180 0.8610 0.7680 ;
      RECT 0.7350 0.1460 0.7850 0.5180 ;
      RECT 0.7350 0.7680 0.7850 0.9140 ;
      RECT 0.2790 0.6180 0.7250 0.6680 ;
      RECT 0.2790 0.6680 0.3290 1.1350 ;
      RECT 0.2790 0.4220 0.3290 0.6180 ;
      RECT 2.0870 0.4090 2.8370 0.4590 ;
      RECT 2.7870 0.4590 2.8370 0.8060 ;
      RECT 2.4070 0.8060 2.8370 0.8560 ;
      RECT 2.4070 0.8560 2.4570 1.1660 ;
      RECT 2.0870 1.1660 2.4570 1.2160 ;
      RECT 1.4030 0.7180 2.0930 0.7680 ;
      RECT 1.0390 1.3080 1.2410 1.3580 ;
      RECT 1.0390 1.1660 1.0890 1.3080 ;
      RECT 1.1910 0.4680 1.2410 1.3080 ;
      RECT 1.0230 0.4180 1.2410 0.4680 ;
      RECT 0.6590 1.4280 1.4850 1.4780 ;
      RECT 0.6590 1.4780 0.7090 1.5840 ;
      RECT 1.8580 1.4280 2.0930 1.4780 ;
    LAYER PO ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 1.2770 1.0320 1.3070 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 1.2770 0.0680 1.3070 0.6420 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 2.0370 1.0320 2.0670 1.6060 ;
      RECT 2.0370 0.0680 2.0670 0.7960 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
  END
END LASX1_LVT

MACRO LASX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.496 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9470 0.6660 1.1190 0.8150 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END D

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.4960 0.0300 ;
        RECT 0.5830 0.0300 0.6330 0.4500 ;
        RECT 0.4310 0.0300 0.4810 0.4500 ;
        RECT 3.1670 0.0300 3.2170 0.2200 ;
        RECT 2.5590 0.0300 2.6090 0.2200 ;
        RECT 2.8630 0.0300 2.9130 0.2200 ;
        RECT 2.4070 0.0300 2.4570 0.2880 ;
        RECT 0.8870 0.2880 2.4570 0.3380 ;
        RECT 0.8870 0.3380 0.9370 0.4620 ;
    END
  END VSS

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.7110 1.1190 2.7610 1.5460 ;
        RECT 2.7110 1.0690 3.2570 1.1190 ;
        RECT 3.1370 1.0090 3.2570 1.0690 ;
        RECT 3.2070 0.4430 3.2570 1.0090 ;
        RECT 2.7110 0.3930 3.2570 0.4430 ;
        RECT 2.7110 0.1480 2.7610 0.3930 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.4960 1.7020 ;
        RECT 2.5590 1.1700 2.6090 1.6420 ;
        RECT 2.8630 1.1700 2.9130 1.6420 ;
        RECT 3.1670 1.3630 3.2170 1.6420 ;
        RECT 0.5590 1.1270 0.6090 1.6420 ;
        RECT 2.4230 1.3780 2.4730 1.6420 ;
        RECT 0.4310 1.0770 0.9370 1.1270 ;
        RECT 1.9760 1.3280 2.4730 1.3780 ;
        RECT 0.4310 0.8610 0.4810 1.0770 ;
        RECT 0.5830 0.8740 0.6330 1.0770 ;
        RECT 0.8870 1.1270 0.9370 1.3430 ;
        RECT 1.9760 1.3150 2.0260 1.3280 ;
        RECT 1.6310 1.2650 2.0260 1.3150 ;
    END
  END VDD

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6170 1.4650 1.7710 1.5750 ;
    END
    ANTENNAGATEAREA 0.018 ;
  END SETB

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9990 0.2920 3.3990 0.3420 ;
        RECT 3.3490 0.3420 3.3990 1.1610 ;
        RECT 3.2890 1.1610 3.4000 1.2210 ;
        RECT 3.0150 1.2210 3.4000 1.2710 ;
        RECT 3.0150 1.2710 3.0650 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 1.3130 0.4050 1.4230 ;
        RECT 0.3550 1.4230 0.4050 1.5840 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  OBS
    LAYER NWELL ;
      RECT 0.2280 0.6770 0.8590 0.6790 ;
      RECT -0.1150 0.6790 3.6110 1.7730 ;
    LAYER M1 ;
      RECT 1.7990 0.6040 2.8530 0.6540 ;
      RECT 1.7990 0.5100 1.8490 0.6040 ;
      RECT 2.1430 0.6540 2.1930 1.0650 ;
      RECT 1.4790 1.0650 2.1930 1.1150 ;
      RECT 1.5550 0.6180 1.6960 0.6680 ;
      RECT 1.6460 0.4600 1.6960 0.6180 ;
      RECT 1.3430 0.4100 2.0170 0.4600 ;
      RECT 1.3430 0.4600 1.3930 0.6060 ;
      RECT 1.3030 0.6060 1.3930 0.6560 ;
      RECT 1.3030 0.6560 1.3530 1.1650 ;
      RECT 1.3030 1.1650 2.0220 1.2150 ;
      RECT 0.7350 0.0960 1.9720 0.1460 ;
      RECT 0.7350 0.5180 0.8610 0.5680 ;
      RECT 0.8110 0.5680 0.8610 0.7180 ;
      RECT 0.7350 0.7180 0.8610 0.7680 ;
      RECT 0.7350 0.1460 0.7850 0.5180 ;
      RECT 0.7350 0.7680 0.7850 0.9140 ;
      RECT 0.2790 0.6180 0.7250 0.6680 ;
      RECT 0.2790 0.6680 0.3290 1.1350 ;
      RECT 0.2790 0.4220 0.3290 0.6180 ;
      RECT 2.9390 0.6040 3.1570 0.6540 ;
      RECT 2.9390 0.6540 2.9890 0.8060 ;
      RECT 2.9390 0.5430 2.9890 0.6040 ;
      RECT 2.4070 0.8060 2.9890 0.8560 ;
      RECT 2.0870 0.4930 2.9890 0.5430 ;
      RECT 2.4070 0.8560 2.4570 1.1660 ;
      RECT 2.0870 1.1660 2.4570 1.2160 ;
      RECT 1.4030 0.7180 2.0930 0.7680 ;
      RECT 1.0390 1.3080 1.2410 1.3580 ;
      RECT 1.0390 1.1660 1.0890 1.3080 ;
      RECT 1.1910 0.4680 1.2410 1.3080 ;
      RECT 1.0230 0.4180 1.2410 0.4680 ;
      RECT 0.6590 1.4280 1.4850 1.4780 ;
      RECT 0.6590 1.4780 0.7090 1.5840 ;
      RECT 1.8580 1.4280 2.0930 1.4780 ;
    LAYER PO ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 1.2770 1.0320 1.3070 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 1.2770 0.0680 1.3070 0.6420 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 2.0370 1.0320 2.0670 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 2.0370 0.0680 2.0670 0.7960 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
  END
END LASX2_LVT

MACRO LATCHX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.04 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9470 0.6660 1.1190 0.8150 ;
    END
    ANTENNAGATEAREA 0.0312 ;
  END D

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.0400 0.0300 ;
        RECT 2.5590 0.0300 2.6090 0.2200 ;
        RECT 0.5830 0.0300 0.6330 0.4500 ;
        RECT 0.4310 0.0300 0.4810 0.4500 ;
        RECT 2.2550 0.0300 2.3050 0.3040 ;
        RECT 0.8870 0.3040 2.3050 0.3540 ;
        RECT 0.8870 0.3540 0.9370 0.4780 ;
    END
  END VSS

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4070 1.0690 2.7910 1.1190 ;
        RECT 2.6810 1.0090 2.7910 1.0690 ;
        RECT 2.4070 1.1190 2.4570 1.5460 ;
        RECT 2.7410 0.3590 2.7910 1.0090 ;
        RECT 2.4070 0.3090 2.7910 0.3590 ;
        RECT 2.4070 0.1480 2.4570 0.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.0400 1.7020 ;
        RECT 2.5590 1.1700 2.6090 1.6420 ;
        RECT 2.2550 1.0840 2.3050 1.6420 ;
        RECT 0.5430 1.1270 0.5930 1.6420 ;
        RECT 1.6620 1.4710 1.7120 1.6420 ;
        RECT 0.4310 1.0770 0.9370 1.1270 ;
        RECT 1.4950 1.4210 1.7120 1.4710 ;
        RECT 0.4310 0.8610 0.4810 1.0770 ;
        RECT 0.5830 0.8740 0.6330 1.0770 ;
        RECT 0.8870 1.1270 0.9370 1.3430 ;
        RECT 1.4950 1.1920 1.5450 1.4210 ;
    END
  END VDD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8330 1.1610 2.9440 1.2210 ;
        RECT 2.7110 1.2210 2.9440 1.2710 ;
        RECT 2.8930 0.2040 2.9430 1.1610 ;
        RECT 2.7110 1.2710 2.7610 1.5460 ;
        RECT 2.6950 0.1540 2.9430 0.2040 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 1.3130 0.4050 1.4230 ;
        RECT 0.3550 1.4230 0.4050 1.5840 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 3.1550 1.7730 ;
      RECT 0.2170 0.6680 0.5420 0.6790 ;
    LAYER M1 ;
      RECT 2.1630 0.6600 2.5490 0.7100 ;
      RECT 2.2530 0.7100 2.3030 0.9080 ;
      RECT 1.6310 0.9080 2.3030 0.9580 ;
      RECT 1.6890 0.5680 1.7390 0.9080 ;
      RECT 1.6310 0.5180 1.7390 0.5680 ;
      RECT 1.3430 0.4100 2.6850 0.4600 ;
      RECT 2.6350 0.4600 2.6850 0.6700 ;
      RECT 1.3430 0.4600 1.3930 1.0280 ;
      RECT 1.4980 0.4600 1.5480 0.6180 ;
      RECT 1.3430 1.0280 1.8490 1.0780 ;
      RECT 1.4980 0.6180 1.6390 0.6680 ;
      RECT 1.7990 1.0780 1.8490 1.2020 ;
      RECT 0.7350 0.0960 2.0930 0.1460 ;
      RECT 0.7350 0.1460 0.7850 0.5180 ;
      RECT 0.7350 0.5180 0.8250 0.5680 ;
      RECT 0.7750 0.5680 0.8250 0.7180 ;
      RECT 0.7350 0.7180 0.8250 0.7680 ;
      RECT 0.7350 0.7680 0.7850 0.9140 ;
      RECT 0.2790 0.6180 0.7250 0.6680 ;
      RECT 0.2790 0.6680 0.3290 1.1350 ;
      RECT 0.2790 0.2250 0.3290 0.6180 ;
      RECT 1.0390 1.3080 1.2410 1.3580 ;
      RECT 1.0390 1.1660 1.0890 1.3080 ;
      RECT 1.1910 0.4680 1.2410 1.3080 ;
      RECT 1.0230 0.4180 1.2410 0.4680 ;
      RECT 0.6430 1.5260 1.4850 1.5760 ;
      RECT 1.9350 0.8080 2.1820 0.8580 ;
      RECT 1.9350 0.5750 1.9850 0.8080 ;
      RECT 1.9350 0.5250 2.1690 0.5750 ;
      RECT 1.4030 0.1960 1.9410 0.2460 ;
      RECT 1.8580 1.5260 2.0930 1.5760 ;
    LAYER PO ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 1.2770 0.0680 1.3070 0.6420 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 1.2770 0.7420 1.3070 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 1.8850 0.7420 1.9150 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 1.8850 0.0680 1.9150 0.6420 ;
  END
END LATCHX1_LVT

MACRO LATCHX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.344 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9470 0.6660 1.1190 0.8150 ;
    END
    ANTENNAGATEAREA 0.0312 ;
  END D

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.3440 0.0300 ;
        RECT 0.5830 0.0300 0.6330 0.4500 ;
        RECT 0.4310 0.0300 0.4810 0.4500 ;
        RECT 3.0150 0.0300 3.0650 0.2200 ;
        RECT 2.7110 0.0300 2.7610 0.2200 ;
        RECT 2.4070 0.0300 2.4570 0.2200 ;
        RECT 2.2550 0.0300 2.3050 0.3040 ;
        RECT 0.8870 0.3040 2.3050 0.3540 ;
        RECT 0.8870 0.3540 0.9370 0.4780 ;
    END
  END VSS

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8330 1.0590 2.9430 1.1190 ;
        RECT 2.5590 1.0090 3.1050 1.0590 ;
        RECT 2.5590 1.0590 2.6090 1.5460 ;
        RECT 3.0550 0.5100 3.1050 1.0090 ;
        RECT 2.5590 0.4600 3.1050 0.5100 ;
        RECT 2.5590 0.1480 2.6090 0.4600 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.3440 1.7020 ;
        RECT 2.2550 1.0840 2.3050 1.6420 ;
        RECT 3.0150 1.3620 3.0650 1.6420 ;
        RECT 2.4070 1.1700 2.4570 1.6420 ;
        RECT 2.7110 1.1700 2.7610 1.6420 ;
        RECT 1.6620 1.4710 1.7120 1.6420 ;
        RECT 0.5430 1.1270 0.5930 1.6420 ;
        RECT 1.4950 1.4210 1.7120 1.4710 ;
        RECT 0.4310 1.0770 0.9370 1.1270 ;
        RECT 1.4950 1.1920 1.5450 1.4210 ;
        RECT 0.4310 0.8610 0.4810 1.0770 ;
        RECT 0.5830 0.8740 0.6330 1.0770 ;
        RECT 0.8870 1.1270 0.9370 1.3430 ;
    END
  END VDD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9850 1.1610 3.0960 1.2210 ;
        RECT 2.8630 1.2210 3.2690 1.2710 ;
        RECT 2.8630 1.2710 2.9130 1.5460 ;
        RECT 3.2190 0.4020 3.2690 1.2210 ;
        RECT 2.8470 0.3520 3.2690 0.4020 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 1.3130 0.4050 1.4230 ;
        RECT 0.3550 1.4230 0.4050 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  OBS
    LAYER NWELL ;
      RECT 0.2280 0.6690 0.5320 0.6790 ;
      RECT -0.1150 0.6790 3.4590 1.7730 ;
    LAYER M1 ;
      RECT 2.3750 0.6040 3.0050 0.6100 ;
      RECT 2.7710 0.6100 3.0050 0.6540 ;
      RECT 1.3430 0.4600 1.3930 1.0280 ;
      RECT 1.4980 0.4600 1.5480 0.6180 ;
      RECT 1.3430 1.0280 1.8490 1.0780 ;
      RECT 1.4980 0.6180 1.6390 0.6680 ;
      RECT 1.7990 1.0780 1.8490 1.2020 ;
      RECT 2.3750 0.4600 2.4250 0.5600 ;
      RECT 1.3430 0.4100 2.4250 0.4600 ;
      RECT 2.3750 0.5600 2.8210 0.6040 ;
      RECT 2.1630 0.6600 2.7010 0.7100 ;
      RECT 2.2530 0.7100 2.3030 0.9080 ;
      RECT 1.6310 0.9080 2.3030 0.9580 ;
      RECT 1.6890 0.5680 1.7390 0.9080 ;
      RECT 1.6310 0.5180 1.7390 0.5680 ;
      RECT 0.7350 0.0960 2.0930 0.1460 ;
      RECT 0.7350 0.1460 0.7850 0.5180 ;
      RECT 0.7350 0.5180 0.8250 0.5680 ;
      RECT 0.7750 0.5680 0.8250 0.7180 ;
      RECT 0.7350 0.7180 0.8250 0.7680 ;
      RECT 0.7350 0.7680 0.7850 0.9140 ;
      RECT 0.2790 0.6180 0.7250 0.6680 ;
      RECT 0.2790 0.6680 0.3290 1.1350 ;
      RECT 0.2790 0.2250 0.3290 0.6180 ;
      RECT 1.0390 1.3080 1.2410 1.3580 ;
      RECT 1.0390 1.1660 1.0890 1.3080 ;
      RECT 1.1910 0.4680 1.2410 1.3080 ;
      RECT 1.0230 0.4180 1.2410 0.4680 ;
      RECT 0.6430 1.5260 1.4850 1.5760 ;
      RECT 1.9350 0.8080 2.1820 0.8580 ;
      RECT 1.9350 0.5750 1.9850 0.8080 ;
      RECT 1.9350 0.5250 2.1690 0.5750 ;
      RECT 1.4030 0.1960 1.9410 0.2460 ;
      RECT 1.8580 1.5260 2.0930 1.5760 ;
    LAYER PO ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 1.2770 0.0680 1.3070 0.6420 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 1.2770 0.7420 1.3070 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 1.8850 0.7420 1.9150 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 1.8850 0.0680 1.9150 0.6420 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
  END
END LATCHX2_LVT

MACRO LNANDX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.368 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0390 0.1060 1.0890 0.5530 ;
        RECT 1.0090 0.5530 1.1290 0.6630 ;
        RECT 1.0790 0.6630 1.1290 1.0170 ;
        RECT 0.4910 1.0170 1.1290 1.0670 ;
        RECT 1.0390 1.0670 1.0890 1.5510 ;
        RECT 0.7350 1.0670 0.7850 1.5510 ;
    END
    ANTENNADIFFAREA 0.086 ;
  END QN

  PIN RIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7950 0.8870 0.9680 0.9370 ;
        RECT 0.8570 0.9370 0.9680 0.9670 ;
        RECT 0.8570 0.8570 0.9680 0.8870 ;
    END
    ANTENNAGATEAREA 0.0216 ;
  END RIN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3880 0.7350 1.0290 0.7850 ;
        RECT 0.5530 0.7850 0.6630 0.8150 ;
        RECT 0.5530 0.7050 0.6630 0.7350 ;
        RECT 0.3880 0.7850 0.4380 1.1230 ;
        RECT 0.5830 0.1060 0.6330 0.7050 ;
        RECT 0.3880 1.1230 0.4810 1.1730 ;
        RECT 0.4310 1.1730 0.4810 1.5510 ;
    END
    ANTENNADIFFAREA 0.0737 ;
  END Q

  PIN SIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.3590 0.5830 ;
        RECT 0.2490 0.5830 0.4210 0.6330 ;
        RECT 0.2490 0.6330 0.3590 0.6630 ;
    END
    ANTENNAGATEAREA 0.0216 ;
  END SIN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.3680 1.7020 ;
        RECT 0.8870 1.2850 0.9370 1.6420 ;
        RECT 0.2790 1.2850 0.3290 1.6420 ;
        RECT 0.5830 1.2850 0.6330 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.3680 0.0300 ;
        RECT 0.7350 0.0300 0.7850 0.4750 ;
        RECT 0.2790 0.0300 0.3290 0.4750 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.0910 0.6790 1.4590 1.7810 ;
    LAYER PO ;
      RECT 1.2770 0.0670 1.3070 1.6010 ;
      RECT 0.9730 0.0670 1.0030 1.6010 ;
      RECT 0.8210 0.0670 0.8510 1.6010 ;
      RECT 1.1250 0.0670 1.1550 1.6010 ;
      RECT 0.6690 0.0670 0.6990 1.6010 ;
      RECT 0.3650 0.0670 0.3950 1.6010 ;
      RECT 0.5170 0.0670 0.5470 1.6010 ;
      RECT 0.2130 0.0670 0.2430 1.6010 ;
      RECT 0.0610 0.0670 0.0910 1.6010 ;
  END
END LNANDX1_LVT

MACRO LNANDX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.976 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN RIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0990 0.8870 1.3330 0.9370 ;
        RECT 1.1610 0.9370 1.2710 0.9670 ;
        RECT 1.1610 0.8570 1.2710 0.8870 ;
    END
    ANTENNAGATEAREA 0.0432 ;
  END RIN

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6170 0.8570 1.7520 0.9670 ;
        RECT 1.7020 0.7880 1.7520 0.8570 ;
        RECT 1.7020 0.9670 1.7520 1.0790 ;
        RECT 0.6430 0.7380 1.7520 0.7880 ;
        RECT 1.0390 1.0790 1.7520 1.1290 ;
        RECT 1.7020 0.5020 1.7520 0.7380 ;
        RECT 1.0390 1.1290 1.0890 1.5670 ;
        RECT 1.6470 1.1290 1.6970 1.5670 ;
        RECT 1.3430 1.1290 1.3930 1.5670 ;
        RECT 1.4950 0.4520 1.7520 0.5020 ;
        RECT 1.4950 0.5020 1.5450 0.5440 ;
    END
    ANTENNADIFFAREA 0.1253 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2390 0.8150 0.2890 1.0790 ;
        RECT 0.2390 1.0790 0.7850 1.1290 ;
        RECT 0.2390 0.7050 0.3590 0.8150 ;
        RECT 0.4310 1.1290 0.4810 1.5670 ;
        RECT 0.7350 1.1290 0.7850 1.5670 ;
        RECT 0.2390 0.6550 0.2890 0.7050 ;
        RECT 0.2390 0.6050 1.6370 0.6550 ;
        RECT 0.7350 0.6550 0.7850 0.6630 ;
        RECT 0.7350 0.4620 0.7850 0.6050 ;
    END
    ANTENNADIFFAREA 0.113 ;
  END Q

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.9760 0.0300 ;
        RECT 1.1910 0.0300 1.2410 0.4020 ;
        RECT 0.4310 0.0300 0.4810 0.4020 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.9760 1.7020 ;
        RECT 1.4950 1.2860 1.5450 1.6420 ;
        RECT 1.1910 1.2860 1.2410 1.6420 ;
        RECT 0.8870 1.2860 0.9370 1.6420 ;
        RECT 0.2790 1.2860 0.3290 1.6420 ;
        RECT 0.5830 1.2860 0.6330 1.6420 ;
    END
  END VDD

  PIN SIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.8870 0.5730 0.9370 ;
        RECT 0.4010 0.9370 0.5110 0.9670 ;
        RECT 0.4010 0.8570 0.5110 0.8870 ;
    END
    ANTENNAGATEAREA 0.0432 ;
  END SIN
  OBS
    LAYER NWELL ;
      RECT -0.0910 0.6790 2.0670 1.7800 ;
    LAYER M1 ;
      RECT 1.3430 0.1860 1.6970 0.2360 ;
      RECT 1.6470 0.2360 1.6970 0.4020 ;
      RECT 1.3430 0.2360 1.3930 0.5050 ;
      RECT 1.0390 0.5050 1.3930 0.5550 ;
      RECT 1.0390 0.1060 1.0890 0.5050 ;
      RECT 0.8870 0.2360 0.9370 0.4020 ;
      RECT 0.5830 0.1860 0.9370 0.2360 ;
      RECT 0.5830 0.2360 0.6330 0.5050 ;
      RECT 0.2790 0.5050 0.6330 0.5550 ;
      RECT 0.2790 0.1060 0.3290 0.5050 ;
    LAYER PO ;
      RECT 1.8850 0.0710 1.9150 1.6030 ;
      RECT 1.4290 0.0710 1.4590 1.6020 ;
      RECT 1.1250 0.0710 1.1550 1.6030 ;
      RECT 1.2770 0.0710 1.3070 1.6020 ;
      RECT 1.5810 0.0710 1.6110 1.6020 ;
      RECT 1.7330 0.0710 1.7630 1.6020 ;
      RECT 0.9730 0.0710 1.0030 1.6020 ;
      RECT 0.0610 0.0710 0.0910 1.6020 ;
      RECT 0.8210 0.0710 0.8510 1.6020 ;
      RECT 0.2130 0.0710 0.2430 1.6020 ;
      RECT 0.5170 0.0710 0.5470 1.6020 ;
      RECT 0.3650 0.0710 0.3950 1.6020 ;
      RECT 0.6690 0.0710 0.6990 1.6020 ;
  END
END LNANDX2_LVT

MACRO LSDNENCLSSX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.368 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6140 0.6490 0.8150 0.7050 ;
        RECT 0.7050 0.7050 0.8150 0.8150 ;
    END
    ANTENNAGATEAREA 0.0366 ;
  END EN

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1900 0.5110 0.2460 0.6520 ;
        RECT 0.0970 0.4010 0.2460 0.5110 ;
        RECT 0.1900 0.6520 0.4230 0.7080 ;
    END
    ANTENNAGATEAREA 0.0366 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0370 0.8820 1.0930 1.5120 ;
        RECT 1.0370 0.8260 1.2710 0.8820 ;
        RECT 1.1540 0.8820 1.2710 0.9670 ;
        RECT 1.1470 0.5720 1.2030 0.8260 ;
        RECT 0.7310 0.5280 1.2030 0.5720 ;
        RECT 0.7310 0.5160 1.1750 0.5280 ;
        RECT 0.7310 0.1260 0.7870 0.5160 ;
        RECT 1.0350 0.1610 1.0910 0.5160 ;
    END
    ANTENNADIFFAREA 0.1672 ;
  END Y

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.3680 0.0300 ;
        RECT 0.5800 0.0300 0.6360 0.2690 ;
        RECT 0.8840 0.0300 0.9400 0.4180 ;
        RECT 0.2760 0.0300 0.3320 0.2600 ;
    END
  END VSS

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.3680 1.7020 ;
        RECT 0.4280 1.2830 0.4840 1.6420 ;
        RECT 0.5830 1.2580 0.6330 1.6420 ;
    END
  END VDDL
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.4810 1.7730 ;
    LAYER M1 ;
      RECT 0.8820 0.6370 1.0320 0.6930 ;
      RECT 0.8820 0.6930 0.9380 0.8840 ;
      RECT 0.2760 0.8840 0.9380 0.9400 ;
      RECT 0.2760 0.9400 0.3320 1.0310 ;
      RECT 0.2760 0.7710 0.3320 0.8840 ;
      RECT 0.4740 0.5960 0.5300 0.8840 ;
      RECT 0.4280 0.5380 0.5300 0.5960 ;
      RECT 0.4280 0.4480 0.4840 0.5380 ;
      RECT 0.7350 1.2540 0.9370 1.3040 ;
      RECT 0.7350 1.3040 0.7850 1.4690 ;
      RECT 0.8870 1.3040 0.9370 1.4690 ;
    LAYER PO ;
      RECT 0.6690 0.0670 0.6990 1.6210 ;
      RECT 0.0610 0.0670 0.0910 1.6210 ;
      RECT 0.2130 0.0670 0.2430 1.6210 ;
      RECT 0.8210 0.0670 0.8510 1.6210 ;
      RECT 0.5170 0.0670 0.5470 1.6210 ;
      RECT 0.3650 0.0670 0.3950 1.6210 ;
      RECT 1.1250 0.0670 1.1550 1.6070 ;
      RECT 1.2770 0.0670 1.3070 1.6070 ;
      RECT 0.9730 0.0670 1.0030 1.6070 ;
  END
END LSDNENCLSSX1_LVT

MACRO LSDNENCLSSX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.52 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 0.7050 0.8150 0.8160 ;
        RECT 0.6140 0.6490 0.8150 0.7050 ;
    END
    ANTENNAGATEAREA 0.0366 ;
  END EN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7310 0.1260 0.7870 0.5160 ;
        RECT 0.7310 0.5160 1.3220 0.5280 ;
        RECT 1.0350 0.1610 1.0910 0.5160 ;
        RECT 0.7310 0.5280 1.3500 0.5720 ;
        RECT 1.2940 0.5720 1.3500 0.7980 ;
        RECT 1.0360 0.7980 1.4240 0.8540 ;
        RECT 1.3080 0.8540 1.4240 0.9670 ;
        RECT 1.0360 0.8540 1.0920 1.2090 ;
    END
    ANTENNADIFFAREA 0.1916 ;
  END Y

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.5200 0.0300 ;
        RECT 0.5800 0.0300 0.6360 0.2690 ;
        RECT 0.8840 0.0300 0.9400 0.4180 ;
        RECT 0.2760 0.0300 0.3320 0.2600 ;
        RECT 1.1870 0.0300 1.2430 0.3950 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2050 0.4010 0.3590 0.5110 ;
        RECT 0.2050 0.5110 0.2610 0.6520 ;
        RECT 0.2050 0.6520 0.4230 0.7080 ;
    END
    ANTENNAGATEAREA 0.0366 ;
  END A

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.5200 1.7020 ;
        RECT 0.4280 1.2830 0.4840 1.6420 ;
        RECT 0.5830 1.2580 0.6330 1.6420 ;
    END
  END VDDL
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.6330 1.7730 ;
    LAYER M1 ;
      RECT 1.1880 1.3110 1.2440 1.5220 ;
      RECT 0.7350 1.2610 1.2440 1.3110 ;
      RECT 1.1880 0.9310 1.2440 1.2610 ;
      RECT 0.8870 1.3110 0.9370 1.4690 ;
      RECT 0.7350 1.3110 0.7850 1.4690 ;
      RECT 0.8820 0.6370 1.1840 0.6930 ;
      RECT 0.8820 0.6930 0.9380 0.8840 ;
      RECT 0.2760 0.8840 0.9380 0.9400 ;
      RECT 0.2760 0.9400 0.3320 1.0310 ;
      RECT 0.2760 0.7710 0.3320 0.8840 ;
      RECT 0.4740 0.5960 0.5300 0.8840 ;
      RECT 0.4280 0.5380 0.5300 0.5960 ;
      RECT 0.4280 0.4480 0.4840 0.5380 ;
    LAYER PO ;
      RECT 0.6690 0.0670 0.6990 1.6210 ;
      RECT 0.0610 0.0670 0.0910 1.6210 ;
      RECT 0.2130 0.0670 0.2430 1.6210 ;
      RECT 0.8210 0.0670 0.8510 1.6210 ;
      RECT 0.5170 0.0670 0.5470 1.6210 ;
      RECT 0.3650 0.0670 0.3950 1.6210 ;
      RECT 1.1250 0.0670 1.1550 1.6070 ;
      RECT 1.2770 0.0670 1.3070 1.6070 ;
      RECT 0.9730 0.0670 1.0030 1.6070 ;
      RECT 1.4290 0.0670 1.4590 1.6070 ;
  END
END LSDNENCLSSX2_LVT

MACRO LSDNENCLSSX4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.824 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0360 0.7980 1.7100 0.8540 ;
        RECT 1.6170 0.8540 1.7270 0.9670 ;
        RECT 1.3400 0.8540 1.3960 1.2090 ;
        RECT 1.0360 0.8540 1.0920 1.2090 ;
        RECT 1.6540 0.7340 1.7100 0.7980 ;
        RECT 1.6530 0.7310 1.7100 0.7340 ;
        RECT 1.6530 0.5720 1.7090 0.7310 ;
        RECT 0.7310 0.5160 1.7090 0.5720 ;
        RECT 0.7310 0.1260 0.7870 0.5160 ;
        RECT 1.0350 0.1610 1.0910 0.5160 ;
        RECT 1.3400 0.1610 1.3960 0.5160 ;
    END
    ANTENNADIFFAREA 0.3404 ;
  END Y

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 0.7050 0.8150 0.8160 ;
        RECT 0.6140 0.6490 0.8150 0.7050 ;
    END
    ANTENNAGATEAREA 0.0366 ;
  END EN

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2070 0.4010 0.3590 0.5110 ;
        RECT 0.2070 0.5110 0.2630 0.6520 ;
        RECT 0.2070 0.6520 0.4230 0.7080 ;
    END
    ANTENNAGATEAREA 0.0366 ;
  END A

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.8240 0.0300 ;
        RECT 0.5800 0.0300 0.6360 0.2690 ;
        RECT 0.8840 0.0300 0.9400 0.4180 ;
        RECT 0.2760 0.0300 0.3320 0.2600 ;
        RECT 1.1870 0.0300 1.2430 0.3950 ;
        RECT 1.4920 0.0300 1.5480 0.3950 ;
    END
  END VSS

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.8240 1.7020 ;
        RECT 0.4280 1.2830 0.4840 1.6420 ;
        RECT 0.5830 1.2580 0.6330 1.6420 ;
    END
  END VDDL
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.9370 1.7730 ;
    LAYER M1 ;
      RECT 1.4920 1.3490 1.5480 1.5220 ;
      RECT 0.8870 1.3040 1.5480 1.3490 ;
      RECT 0.7350 1.2990 1.5480 1.3040 ;
      RECT 1.4920 1.1980 1.5480 1.2990 ;
      RECT 0.8870 1.3490 0.9370 1.4690 ;
      RECT 0.7350 1.3040 0.7850 1.4690 ;
      RECT 0.7350 1.2540 0.9370 1.2990 ;
      RECT 1.1880 1.3490 1.2440 1.5220 ;
      RECT 1.1880 1.1960 1.2440 1.2990 ;
      RECT 0.8820 0.6370 1.5000 0.6930 ;
      RECT 0.8820 0.6930 0.9380 0.8840 ;
      RECT 0.2760 0.8840 0.9380 0.9400 ;
      RECT 0.2760 0.9400 0.3320 1.0310 ;
      RECT 0.2760 0.7710 0.3320 0.8840 ;
      RECT 0.4740 0.5960 0.5300 0.8840 ;
      RECT 0.4280 0.5380 0.5300 0.5960 ;
      RECT 0.4280 0.4480 0.4840 0.5380 ;
    LAYER PO ;
      RECT 1.5810 0.0670 1.6110 1.6070 ;
      RECT 0.6690 0.0670 0.6990 1.6210 ;
      RECT 0.0610 0.0670 0.0910 1.6210 ;
      RECT 0.2130 0.0670 0.2430 1.6210 ;
      RECT 0.8210 0.0670 0.8510 1.6210 ;
      RECT 0.5170 0.0670 0.5470 1.6210 ;
      RECT 0.3650 0.0670 0.3950 1.6210 ;
      RECT 1.1250 0.0670 1.1550 1.6070 ;
      RECT 1.2770 0.0670 1.3070 1.6070 ;
      RECT 0.9730 0.0670 1.0030 1.6070 ;
      RECT 1.7330 0.0670 1.7630 1.6070 ;
      RECT 1.4290 0.0670 1.4590 1.6070 ;
  END
END LSDNENCLSSX4_LVT

MACRO LSDNENCLSSX8_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.432 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7310 0.5160 2.2690 0.5720 ;
        RECT 0.7310 0.1260 0.7870 0.5160 ;
        RECT 2.2130 0.5720 2.2690 0.7310 ;
        RECT 1.9480 0.1610 2.0040 0.5160 ;
        RECT 1.6440 0.1610 1.7000 0.5160 ;
        RECT 1.0350 0.1610 1.0910 0.5160 ;
        RECT 1.3400 0.1610 1.3960 0.5160 ;
        RECT 2.2130 0.7310 2.2700 0.7340 ;
        RECT 2.2140 0.7340 2.2700 0.7980 ;
        RECT 1.0360 0.7980 2.2700 0.8070 ;
        RECT 1.0360 0.8070 2.3350 0.8540 ;
        RECT 2.2150 0.8540 2.3350 0.9670 ;
        RECT 1.6440 0.8540 1.7000 1.2090 ;
        RECT 1.9480 0.8540 2.0040 1.2090 ;
        RECT 1.3400 0.8540 1.3960 1.2090 ;
        RECT 1.0360 0.8540 1.0920 1.2090 ;
    END
    ANTENNADIFFAREA 0.638 ;
  END Y

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6140 0.6490 0.8150 0.7050 ;
        RECT 0.7050 0.7050 0.8150 0.8150 ;
    END
    ANTENNAGATEAREA 0.0366 ;
  END EN

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2130 0.5110 0.2690 0.6510 ;
        RECT 0.2130 0.4010 0.3590 0.5110 ;
        RECT 0.2130 0.6510 0.3320 0.6520 ;
        RECT 0.2130 0.6520 0.4230 0.7070 ;
        RECT 0.2970 0.7070 0.4230 0.7080 ;
    END
    ANTENNAGATEAREA 0.0366 ;
  END A

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.4320 0.0300 ;
        RECT 0.5800 0.0300 0.6360 0.2690 ;
        RECT 2.1010 0.0300 2.1570 0.3950 ;
        RECT 0.8840 0.0300 0.9400 0.4180 ;
        RECT 0.2760 0.0300 0.3320 0.2600 ;
        RECT 1.1870 0.0300 1.2430 0.3950 ;
        RECT 1.4920 0.0300 1.5480 0.3950 ;
        RECT 1.7960 0.0300 1.8520 0.3950 ;
    END
  END VSS

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.4320 1.7020 ;
        RECT 0.4280 1.2830 0.4840 1.6420 ;
        RECT 0.5830 1.2580 0.6330 1.6420 ;
    END
  END VDDL
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 2.5450 1.7730 ;
    LAYER M1 ;
      RECT 2.1000 1.3490 2.1560 1.5220 ;
      RECT 0.8870 1.3040 2.1560 1.3490 ;
      RECT 0.7350 1.2990 2.1560 1.3040 ;
      RECT 2.1000 1.1980 2.1560 1.2990 ;
      RECT 0.8870 1.3490 0.9370 1.4690 ;
      RECT 0.7350 1.3040 0.7850 1.4690 ;
      RECT 0.7350 1.2540 0.9370 1.2990 ;
      RECT 1.1880 1.3490 1.2440 1.5220 ;
      RECT 1.1880 1.1960 1.2440 1.2990 ;
      RECT 1.4920 1.3490 1.5480 1.5220 ;
      RECT 1.4920 1.1980 1.5480 1.2990 ;
      RECT 1.7960 1.3490 1.8520 1.5220 ;
      RECT 1.7960 1.1960 1.8520 1.2990 ;
      RECT 0.8820 0.6370 2.1070 0.6930 ;
      RECT 0.8820 0.6930 0.9380 0.8840 ;
      RECT 0.2760 0.8840 0.9380 0.9400 ;
      RECT 0.2760 0.9400 0.3320 1.0310 ;
      RECT 0.2760 0.7710 0.3320 0.8840 ;
      RECT 0.4740 0.5960 0.5300 0.8840 ;
      RECT 0.4280 0.5380 0.5300 0.5960 ;
      RECT 0.4280 0.4480 0.4840 0.5380 ;
    LAYER PO ;
      RECT 2.3410 0.0670 2.3710 1.6070 ;
      RECT 1.5810 0.0670 1.6110 1.6070 ;
      RECT 0.6690 0.0670 0.6990 1.6210 ;
      RECT 0.0610 0.0670 0.0910 1.6210 ;
      RECT 0.2130 0.0670 0.2430 1.6210 ;
      RECT 0.8210 0.0670 0.8510 1.6210 ;
      RECT 0.5170 0.0670 0.5470 1.6210 ;
      RECT 0.3650 0.0670 0.3950 1.6210 ;
      RECT 1.1250 0.0670 1.1550 1.6070 ;
      RECT 1.2770 0.0670 1.3070 1.6070 ;
      RECT 0.9730 0.0670 1.0030 1.6070 ;
      RECT 1.7330 0.0670 1.7630 1.6070 ;
      RECT 2.1890 0.0670 2.2190 1.6070 ;
      RECT 2.0370 0.0670 2.0670 1.6070 ;
      RECT 1.8850 0.0670 1.9150 1.6070 ;
      RECT 1.4290 0.0670 1.4590 1.6070 ;
  END
END LSDNENCLSSX8_LVT

MACRO LSDNENCLX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.128 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9420 1.1470 1.1330 1.2810 ;
    END
    ANTENNAGATEAREA 0.048 ;
  END EN

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.1280 0.0300 ;
        RECT 1.7990 0.0300 1.8490 0.4850 ;
        RECT 1.0390 0.0300 1.0890 0.5050 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 2.1280 3.3740 ;
    END
  END VDDL

  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 3.0100 2.1280 3.0700 ;
        RECT 1.1620 3.0700 1.2720 3.1440 ;
        RECT 1.1620 2.9360 1.2720 3.0100 ;
        RECT 0.8870 2.5250 0.9370 3.0100 ;
        RECT 1.1910 2.5200 1.2410 2.9360 ;
    END
  END VDDH

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.1280 1.7020 ;
        RECT 1.0390 1.4960 1.0890 1.6420 ;
        RECT 1.0390 1.7020 1.0890 2.1290 ;
        RECT 0.5830 1.4850 0.6330 1.6420 ;
        RECT 1.7990 1.3030 1.8490 1.6420 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7850 0.8310 0.8350 0.8420 ;
        RECT 0.7850 0.8420 0.9870 0.9760 ;
        RECT 0.4310 0.7810 0.8350 0.8310 ;
        RECT 0.7850 0.9760 0.8350 1.1980 ;
        RECT 0.4310 0.2280 0.4810 0.7810 ;
        RECT 0.7350 0.2300 0.7850 0.7810 ;
        RECT 0.7350 1.1980 0.8350 1.2620 ;
        RECT 0.7350 1.2620 0.7850 1.5230 ;
        RECT 0.7350 1.5230 0.9370 1.5730 ;
        RECT 0.8870 1.4780 0.9370 1.5230 ;
    END
    ANTENNADIFFAREA 0.1734 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7940 2.2130 1.1600 2.2630 ;
        RECT 0.9970 2.2630 1.1600 2.3650 ;
    END
    ANTENNAGATEAREA 0.0261 ;
  END A
  OBS
    LAYER NWELL ;
      RECT -0.1150 3.2240 2.2430 3.4590 ;
      RECT -0.1150 2.3510 0.1150 3.2240 ;
      RECT 2.0130 2.3510 2.2430 3.2240 ;
      RECT 0.5750 2.2340 1.4250 2.7640 ;
      RECT -0.1150 -0.1150 2.2430 0.9930 ;
    LAYER M1 ;
      RECT 0.8870 0.6640 1.2410 0.7140 ;
      RECT 1.1910 0.2300 1.2410 0.6640 ;
      RECT 0.8870 0.1380 0.9370 0.6640 ;
      RECT 0.5830 0.0880 0.9370 0.1380 ;
      RECT 0.5830 0.1380 0.6330 0.6310 ;
      RECT 0.9470 1.0280 1.1810 1.0780 ;
      RECT 0.6750 2.4230 1.0890 2.4730 ;
      RECT 1.0390 2.4730 1.0890 2.6900 ;
      RECT 0.6750 2.2630 0.7250 2.4230 ;
      RECT 0.4900 2.2130 0.7250 2.2630 ;
      RECT 0.6750 2.1280 0.7250 2.2130 ;
      RECT 0.6750 2.0780 0.9370 2.1280 ;
      RECT 0.8870 1.9760 0.9370 2.0780 ;
      RECT 0.7350 2.4730 0.7850 2.6900 ;
      RECT 0.4910 1.0280 0.7250 1.0780 ;
    LAYER PO ;
      RECT 1.7330 0.0690 1.7630 2.7800 ;
      RECT 0.3650 0.0890 0.3950 2.7800 ;
      RECT 1.1250 0.0870 1.1550 2.7780 ;
      RECT 1.8850 0.0690 1.9150 2.7800 ;
      RECT 0.8210 1.7710 0.8510 2.7820 ;
      RECT 0.9730 0.0890 1.0030 1.6690 ;
      RECT 1.5810 0.0690 1.6110 2.7800 ;
      RECT 1.2770 0.0750 1.3070 2.7800 ;
      RECT 1.4290 0.0750 1.4590 2.7800 ;
      RECT 2.0370 0.0740 2.0670 2.7800 ;
      RECT 0.9730 1.7690 1.0030 2.7820 ;
      RECT 0.8210 0.0780 0.8510 1.6700 ;
      RECT 0.0610 0.0890 0.0910 2.7800 ;
      RECT 0.6690 0.0890 0.6990 2.7810 ;
      RECT 0.5170 0.0890 0.5470 2.7800 ;
      RECT 0.2130 0.0890 0.2430 2.7800 ;
  END
END LSDNENCLX1_LVT

MACRO LSDNENCLX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.28 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.2800 1.7020 ;
        RECT 1.3140 1.7020 1.4240 1.7750 ;
        RECT 1.3140 1.5680 1.4240 1.6420 ;
        RECT 0.8870 1.5170 0.9370 1.6420 ;
        RECT 1.6470 1.3630 1.6970 1.6420 ;
        RECT 0.4310 1.5060 0.4810 1.6420 ;
        RECT 1.9510 1.3150 2.0010 1.6420 ;
        RECT 1.0390 1.7020 1.0890 2.1290 ;
        RECT 1.3430 1.5240 1.3930 1.5680 ;
    END
  END VSS

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7900 1.1200 0.9810 1.2710 ;
    END
    ANTENNAGATEAREA 0.063 ;
  END EN

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.2800 0.0300 ;
        RECT 1.6470 0.0300 1.6970 0.3450 ;
        RECT 0.8870 0.0300 0.9370 0.5050 ;
        RECT 1.3430 0.0300 1.3930 0.3450 ;
        RECT 1.9510 0.0300 2.0010 0.4850 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 2.2800 3.3740 ;
    END
  END VDDL

  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 3.0100 2.2800 3.0700 ;
        RECT 1.3140 3.0700 1.4240 3.1430 ;
        RECT 1.3140 2.9360 1.4240 3.0100 ;
        RECT 1.0390 2.5250 1.0890 3.0100 ;
        RECT 1.3430 2.5200 1.3930 2.9360 ;
    END
  END VDDH

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9080 0.6700 1.9580 0.6940 ;
        RECT 1.9080 0.6940 2.0590 0.8280 ;
        RECT 1.4950 0.6200 1.9580 0.6700 ;
        RECT 1.9080 0.8280 1.9580 1.2010 ;
        RECT 1.7990 0.2170 1.8490 0.6200 ;
        RECT 1.4950 0.1850 1.5450 0.6200 ;
        RECT 1.4950 1.2010 1.9580 1.2510 ;
        RECT 1.7990 1.2510 1.8490 1.5730 ;
        RECT 1.4950 1.2510 1.5450 1.5730 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9460 2.2130 1.3120 2.2630 ;
        RECT 1.1490 2.2630 1.3120 2.3650 ;
    END
    ANTENNAGATEAREA 0.0261 ;
  END A
  OBS
    LAYER NWELL ;
      RECT -0.1150 3.2240 2.3950 3.4590 ;
      RECT -0.1150 2.3510 0.1150 3.2240 ;
      RECT 2.1650 2.3510 2.3950 3.2240 ;
      RECT 0.5750 2.2340 1.6170 2.7640 ;
      RECT -0.1150 -0.1150 2.3950 0.9930 ;
    LAYER M1 ;
      RECT 1.3830 1.0330 1.8200 1.0830 ;
      RECT 1.3830 1.0830 1.4330 1.2010 ;
      RECT 1.3830 0.7050 1.4330 1.0330 ;
      RECT 1.1910 1.2010 1.4330 1.2510 ;
      RECT 1.1720 0.6550 1.4330 0.7050 ;
      RECT 1.1910 1.2510 1.2410 1.3610 ;
      RECT 1.0390 0.2300 1.0890 0.6640 ;
      RECT 0.7350 0.6640 1.0890 0.7140 ;
      RECT 0.7350 0.1470 0.7850 0.6640 ;
      RECT 0.4310 0.0970 0.7850 0.1470 ;
      RECT 0.4310 0.1470 0.4810 0.6310 ;
      RECT 0.8270 2.4230 1.2410 2.4730 ;
      RECT 1.1910 2.4730 1.2410 2.6900 ;
      RECT 0.8270 2.2850 0.8770 2.4230 ;
      RECT 0.7660 2.2630 0.8770 2.2850 ;
      RECT 0.3380 2.2130 0.8770 2.2630 ;
      RECT 0.7660 2.1840 0.8770 2.2130 ;
      RECT 0.8270 2.1280 0.8770 2.1840 ;
      RECT 0.8870 2.4730 0.9370 2.6900 ;
      RECT 0.8270 2.0780 0.9370 2.1280 ;
      RECT 0.8870 1.9760 0.9370 2.0780 ;
      RECT 1.2200 1.0280 1.3330 1.0780 ;
      RECT 0.7350 1.4200 0.7850 1.5840 ;
      RECT 0.2790 0.2280 0.3290 0.7810 ;
      RECT 0.6330 0.8310 0.6830 0.9010 ;
      RECT 0.6330 0.9510 0.6830 1.1980 ;
      RECT 0.2790 0.7810 0.6830 0.8310 ;
      RECT 0.5830 1.1980 0.6830 1.2620 ;
      RECT 0.5830 0.2300 0.6330 0.7810 ;
      RECT 0.5830 1.2620 0.6330 1.3700 ;
      RECT 0.5830 1.4200 0.6330 1.5840 ;
      RECT 0.5830 1.3700 1.0890 1.4200 ;
      RECT 1.0390 1.4200 1.0890 1.5840 ;
      RECT 1.2200 0.9510 1.2700 1.0280 ;
      RECT 0.6330 0.9010 1.2700 0.9510 ;
      RECT 0.7950 1.0010 1.0290 1.0510 ;
      RECT 0.3390 1.0280 0.5730 1.0780 ;
    LAYER PO ;
      RECT 0.6690 0.0780 0.6990 2.7810 ;
      RECT 1.8850 0.0690 1.9150 2.7800 ;
      RECT 0.3650 0.0890 0.3950 2.7800 ;
      RECT 1.1250 0.0870 1.1550 2.7780 ;
      RECT 0.9730 0.0780 1.0030 1.7850 ;
      RECT 2.0370 0.0690 2.0670 2.7800 ;
      RECT 1.5810 0.0660 1.6110 2.7800 ;
      RECT 1.2770 0.0750 1.3070 2.7800 ;
      RECT 1.4290 0.0750 1.4590 2.7800 ;
      RECT 2.1890 0.0740 2.2190 2.7800 ;
      RECT 0.8210 0.0780 0.8510 2.7800 ;
      RECT 1.7330 0.0660 1.7630 2.7800 ;
      RECT 0.2130 0.0890 0.2430 2.7800 ;
      RECT 0.9730 1.9210 1.0030 2.7820 ;
      RECT 0.0610 0.0890 0.0910 2.7800 ;
      RECT 0.5170 0.0890 0.5470 2.7800 ;
  END
END LSDNENCLX2_LVT

MACRO ISOLORAOX4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.408 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.7350 0.5110 0.7850 ;
        RECT 0.4010 0.7850 0.5110 0.8150 ;
        RECT 0.4010 0.7050 0.5110 0.7350 ;
    END
    ANTENNAGATEAREA 0.0186 ;
  END D

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.4080 1.7020 ;
        RECT 0.4310 1.1960 0.4810 1.6420 ;
    END
  END VDD

  PIN ISO
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7070 1.3430 1.9410 1.3930 ;
        RECT 1.7690 1.3930 1.8790 1.4230 ;
        RECT 1.7690 1.3130 1.8790 1.3430 ;
    END
    ANTENNAGATEAREA 0.0318 ;
  END ISO

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.4080 0.0300 ;
        RECT 2.8630 0.0300 2.9130 0.2030 ;
        RECT 3.1670 0.0300 3.2170 0.2030 ;
        RECT 0.4310 0.0300 0.4810 0.2950 ;
        RECT 1.6470 0.0300 1.6970 0.2130 ;
        RECT 2.5590 0.0300 2.6090 0.2030 ;
        RECT 1.9510 0.0300 2.0010 0.2160 ;
        RECT 1.3430 0.0300 1.3930 0.2240 ;
        RECT 2.2550 0.0300 2.3050 0.2030 ;
    END
  END VSS

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4410 0.4010 3.5520 0.4780 ;
        RECT 3.3190 0.4780 3.5520 0.5280 ;
        RECT 3.4610 0.3030 3.5110 0.4010 ;
        RECT 3.3190 0.5280 3.3690 0.6620 ;
        RECT 2.1030 0.2530 3.5110 0.3030 ;
        RECT 2.1030 0.6620 3.3690 0.7120 ;
        RECT 3.3190 0.1790 3.3690 0.2530 ;
        RECT 3.0150 0.1790 3.0650 0.2530 ;
        RECT 2.1030 0.1790 2.1530 0.2530 ;
        RECT 2.7110 0.1790 2.7610 0.2530 ;
        RECT 2.4070 0.1790 2.4570 0.2530 ;
        RECT 3.0150 0.7120 3.0650 1.0280 ;
        RECT 2.4070 0.7120 2.4570 1.0280 ;
        RECT 2.7110 0.7120 2.7610 1.0280 ;
        RECT 2.1030 0.7120 2.1530 1.0280 ;
        RECT 3.3190 0.7120 3.3690 1.0280 ;
    END
    ANTENNADIFFAREA 0.3476 ;
  END Q

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 3.4410 0.7050 3.5510 0.8150 ;
        RECT 3.4710 0.6830 3.5210 0.7050 ;
        RECT 3.4710 0.8150 3.5210 1.0780 ;
        RECT 1.7990 1.0780 3.5210 1.1280 ;
        RECT 1.7990 0.8540 1.8490 1.0780 ;
        RECT 2.8630 0.7620 2.9130 1.0780 ;
        RECT 3.1670 0.7620 3.2170 1.0780 ;
        RECT 2.5590 0.7620 2.6090 1.0780 ;
        RECT 2.2550 0.7620 2.3050 1.0780 ;
    END
  END VDDG
  OBS
    LAYER NWELL ;
      RECT -0.0910 1.5430 4.5230 1.7730 ;
      RECT -0.0910 0.6790 0.7190 1.5430 ;
      RECT 4.2350 0.6790 4.5230 1.5430 ;
      RECT 1.1790 0.4530 3.7750 1.0830 ;
    LAYER M1 ;
      RECT 0.2390 0.9810 0.5730 1.0310 ;
      RECT 0.2390 1.0310 0.2890 1.0960 ;
      RECT 0.2390 0.5040 0.3290 0.5540 ;
      RECT 0.2390 1.0960 0.3290 1.1700 ;
      RECT 0.2790 0.1210 0.3290 0.5040 ;
      RECT 0.2790 1.1700 0.3290 1.5540 ;
      RECT 0.2390 0.5540 0.2890 0.9810 ;
      RECT 0.7950 1.3430 1.6370 1.3930 ;
      RECT 0.7950 0.7480 0.8450 1.3430 ;
      RECT 0.6230 0.6980 0.8450 0.7480 ;
      RECT 0.7950 0.6970 0.8450 0.6980 ;
      RECT 0.6230 0.7480 0.6730 1.1200 ;
      RECT 0.6230 0.5740 0.6730 0.6980 ;
      RECT 0.5830 1.1200 0.6730 1.1700 ;
      RECT 0.5830 0.5240 0.6730 0.5740 ;
      RECT 0.5830 1.1700 0.6330 1.5610 ;
      RECT 0.5830 0.1140 0.6330 0.5240 ;
      RECT 1.6470 0.6700 2.0010 0.7200 ;
      RECT 1.9510 0.7200 2.0010 1.0280 ;
      RECT 1.6470 0.7200 1.6970 1.0780 ;
      RECT 1.3430 1.0780 1.6970 1.1280 ;
      RECT 1.3430 0.7620 1.3930 1.0780 ;
      RECT 1.4950 0.3770 3.3090 0.4270 ;
      RECT 1.4950 0.4270 1.5450 1.0280 ;
      RECT 1.4950 0.1260 1.5450 0.3770 ;
      RECT 1.7990 0.1310 1.8490 0.3770 ;
    LAYER PO ;
      RECT 4.3170 0.0710 4.3470 1.6040 ;
      RECT 1.4290 0.0710 1.4590 1.6040 ;
      RECT 2.4930 0.0710 2.5230 1.6040 ;
      RECT 4.1650 0.0710 4.1950 1.6040 ;
      RECT 1.5810 0.0710 1.6110 1.6040 ;
      RECT 1.8850 0.0710 1.9150 1.6040 ;
      RECT 1.7330 0.0710 1.7630 1.6040 ;
      RECT 2.1890 0.0710 2.2190 1.6040 ;
      RECT 3.1010 0.0710 3.1310 1.6040 ;
      RECT 2.3410 0.0710 2.3710 1.6040 ;
      RECT 2.6450 0.0710 2.6750 1.6040 ;
      RECT 2.7970 0.0710 2.8270 1.6040 ;
      RECT 2.9490 0.0710 2.9790 1.6040 ;
      RECT 0.2130 0.0710 0.2430 1.6040 ;
      RECT 3.5570 0.0710 3.5870 1.6040 ;
      RECT 3.2530 0.0710 3.2830 1.6040 ;
      RECT 3.8610 0.0710 3.8910 1.6040 ;
      RECT 4.0130 0.0710 4.0430 1.6040 ;
      RECT 3.7090 0.0710 3.7390 1.6040 ;
      RECT 3.4050 0.0710 3.4350 1.6040 ;
      RECT 0.0610 0.0710 0.0910 1.6040 ;
      RECT 0.5170 0.0710 0.5470 1.6040 ;
      RECT 0.3650 0.0710 0.3950 1.6040 ;
      RECT 0.6690 0.0710 0.6990 1.6040 ;
      RECT 0.8210 0.0710 0.8510 1.6040 ;
      RECT 2.0370 0.0720 2.0670 1.6040 ;
      RECT 0.9730 0.0710 1.0030 1.6040 ;
      RECT 1.2770 0.0710 1.3070 1.6040 ;
      RECT 1.1250 0.0710 1.1550 1.6040 ;
  END
END ISOLORAOX4_LVT

MACRO ISOLORAOX8_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.928 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.9610 0.4010 5.0720 0.4780 ;
        RECT 4.8390 0.4780 5.0720 0.5280 ;
        RECT 4.9810 0.3030 5.0310 0.4010 ;
        RECT 4.8390 0.5280 4.8890 0.5360 ;
        RECT 2.4070 0.2530 5.0310 0.3030 ;
        RECT 2.4070 0.5360 4.8890 0.5860 ;
        RECT 2.7110 0.1790 2.7610 0.2530 ;
        RECT 2.4070 0.1790 2.4570 0.2530 ;
        RECT 3.3190 0.1790 3.3690 0.2530 ;
        RECT 3.6230 0.1790 3.6730 0.2530 ;
        RECT 3.0150 0.1790 3.0650 0.2530 ;
        RECT 3.9270 0.1790 3.9770 0.2530 ;
        RECT 4.2310 0.1790 4.2810 0.2530 ;
        RECT 4.8390 0.1790 4.8890 0.2530 ;
        RECT 4.5350 0.1790 4.5850 0.2530 ;
        RECT 3.0150 0.5860 3.0650 1.0280 ;
        RECT 2.4070 0.5860 2.4570 1.0280 ;
        RECT 3.6230 0.5860 3.6730 1.0280 ;
        RECT 3.3190 0.5860 3.3690 1.0280 ;
        RECT 2.7110 0.5860 2.7610 1.0280 ;
        RECT 4.5350 0.5860 4.5850 1.0280 ;
        RECT 4.2310 0.5860 4.2810 1.0280 ;
        RECT 3.9270 0.5860 3.9770 1.0280 ;
        RECT 4.8390 0.5860 4.8890 1.0280 ;
    END
    ANTENNADIFFAREA 0.6452 ;
  END Q

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 5.9280 0.0300 ;
        RECT 2.5590 0.0300 2.6090 0.2030 ;
        RECT 0.4310 0.0300 0.4810 0.2950 ;
        RECT 3.4710 0.0300 3.5210 0.2030 ;
        RECT 3.1670 0.0300 3.2170 0.2030 ;
        RECT 2.8630 0.0300 2.9130 0.2030 ;
        RECT 1.6470 0.0300 1.6970 0.2130 ;
        RECT 1.9510 0.0300 2.0010 0.2160 ;
        RECT 1.3430 0.0300 1.3930 0.2240 ;
        RECT 2.2550 0.0300 2.3050 0.2130 ;
        RECT 4.6870 0.0300 4.7370 0.2030 ;
        RECT 4.3830 0.0300 4.4330 0.2030 ;
        RECT 4.0790 0.0300 4.1290 0.2030 ;
        RECT 3.7750 0.0300 3.8250 0.2030 ;
    END
  END VSS

  PIN ISO
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8590 1.3430 2.2450 1.3930 ;
        RECT 1.9210 1.3930 2.0310 1.4230 ;
        RECT 1.9210 1.3130 2.0310 1.3430 ;
    END
    ANTENNAGATEAREA 0.0504 ;
  END ISO

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 5.9280 1.7020 ;
        RECT 0.4310 1.1960 0.4810 1.6420 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.7350 0.5110 0.7850 ;
        RECT 0.4010 0.7850 0.5110 0.8150 ;
        RECT 0.4010 0.7050 0.5110 0.7350 ;
    END
    ANTENNAGATEAREA 0.0186 ;
  END D

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 4.9610 0.7050 5.0710 0.8150 ;
        RECT 4.9910 0.6830 5.0410 0.7050 ;
        RECT 4.9910 0.8150 5.0410 1.0790 ;
        RECT 1.9510 1.0790 5.0410 1.1290 ;
        RECT 2.8630 0.6700 2.9130 1.0790 ;
        RECT 2.5590 0.6700 2.6090 1.0790 ;
        RECT 1.9510 0.6700 2.0010 1.0790 ;
        RECT 3.4710 0.6700 3.5210 1.0790 ;
        RECT 3.1670 0.6700 3.2170 1.0790 ;
        RECT 4.6870 0.6700 4.7370 1.0790 ;
        RECT 2.2550 0.6700 2.3050 1.0790 ;
        RECT 4.3830 0.6700 4.4330 1.0790 ;
        RECT 3.7750 0.6700 3.8250 1.0790 ;
        RECT 4.0790 0.6700 4.1290 1.0790 ;
    END
  END VDDG
  OBS
    LAYER NWELL ;
      RECT 1.1790 0.4530 5.2950 1.0830 ;
      RECT -0.0910 1.5430 6.0420 1.7730 ;
      RECT -0.0910 0.6790 0.7190 1.5430 ;
      RECT 5.7550 0.6790 6.0420 1.5430 ;
    LAYER M1 ;
      RECT 0.7950 1.3430 1.7890 1.3930 ;
      RECT 0.7950 0.7480 0.8450 1.3430 ;
      RECT 0.6230 0.6980 0.8450 0.7480 ;
      RECT 0.7950 0.6970 0.8450 0.6980 ;
      RECT 0.6230 0.5740 0.6730 0.6980 ;
      RECT 0.6230 0.7480 0.6730 1.1200 ;
      RECT 0.5830 0.5240 0.6730 0.5740 ;
      RECT 0.5830 1.1200 0.6730 1.1700 ;
      RECT 0.5830 0.1140 0.6330 0.5240 ;
      RECT 0.5830 1.1700 0.6330 1.5610 ;
      RECT 0.2390 0.9810 0.5730 1.0310 ;
      RECT 0.2390 1.0310 0.2890 1.0960 ;
      RECT 0.2390 0.5040 0.3290 0.5540 ;
      RECT 0.2390 1.0960 0.3290 1.1700 ;
      RECT 0.2790 0.1210 0.3290 0.5040 ;
      RECT 0.2790 1.1700 0.3290 1.5540 ;
      RECT 0.2390 0.5540 0.2890 0.9810 ;
      RECT 1.4950 0.3770 4.8290 0.4270 ;
      RECT 1.4950 0.1260 1.5450 0.3770 ;
      RECT 1.4950 0.4270 1.5450 0.5520 ;
      RECT 1.3430 0.6020 1.3930 1.1070 ;
      RECT 1.7990 0.1310 1.8490 0.3770 ;
      RECT 1.3430 0.5520 1.6970 0.6020 ;
      RECT 1.6470 0.6020 1.6970 1.0280 ;
      RECT 2.1030 0.1260 2.1530 0.3770 ;
      RECT 1.7990 0.5620 2.1530 0.6120 ;
      RECT 2.1030 0.6120 2.1530 1.0290 ;
      RECT 1.7990 0.6120 1.8490 1.0790 ;
      RECT 1.4950 1.0790 1.8490 1.1290 ;
      RECT 1.4950 0.6530 1.5450 1.0790 ;
    LAYER PO ;
      RECT 5.2290 0.0710 5.2590 1.6040 ;
      RECT 5.3810 0.0710 5.4110 1.6040 ;
      RECT 5.5330 0.0710 5.5630 1.6040 ;
      RECT 5.6850 0.0710 5.7150 1.6040 ;
      RECT 5.8370 0.0710 5.8670 1.6040 ;
      RECT 4.7730 0.0710 4.8030 1.6040 ;
      RECT 2.0370 0.0710 2.0670 1.6040 ;
      RECT 2.1890 0.0710 2.2190 1.6040 ;
      RECT 4.9250 0.0710 4.9550 1.6040 ;
      RECT 2.6450 0.0710 2.6750 1.6040 ;
      RECT 3.4050 0.0710 3.4350 1.6040 ;
      RECT 2.4930 0.0710 2.5230 1.6040 ;
      RECT 1.7330 0.0710 1.7630 1.6040 ;
      RECT 1.8850 0.0710 1.9150 1.6040 ;
      RECT 1.5810 0.0710 1.6110 1.6040 ;
      RECT 1.4290 0.0710 1.4590 1.6040 ;
      RECT 2.7970 0.0710 2.8270 1.6040 ;
      RECT 1.1250 0.0710 1.1550 1.6040 ;
      RECT 1.2770 0.0710 1.3070 1.6040 ;
      RECT 0.9730 0.0710 1.0030 1.6040 ;
      RECT 2.3410 0.0720 2.3710 1.6040 ;
      RECT 0.8210 0.0710 0.8510 1.6040 ;
      RECT 0.6690 0.0710 0.6990 1.6040 ;
      RECT 0.3650 0.0710 0.3950 1.6040 ;
      RECT 0.5170 0.0710 0.5470 1.6040 ;
      RECT 0.0610 0.0710 0.0910 1.6040 ;
      RECT 3.7090 0.0710 3.7390 1.6040 ;
      RECT 4.0130 0.0710 4.0430 1.6040 ;
      RECT 4.4690 0.0710 4.4990 1.6040 ;
      RECT 4.6210 0.0710 4.6510 1.6040 ;
      RECT 4.3170 0.0710 4.3470 1.6040 ;
      RECT 4.1650 0.0710 4.1950 1.6040 ;
      RECT 3.5570 0.0710 3.5870 1.6040 ;
      RECT 3.8610 0.0710 3.8910 1.6040 ;
      RECT 0.2130 0.0710 0.2430 1.6040 ;
      RECT 3.2530 0.0710 3.2830 1.6040 ;
      RECT 3.1010 0.0710 3.1310 1.6040 ;
      RECT 2.9490 0.0710 2.9790 1.6040 ;
      RECT 5.0770 0.0710 5.1070 1.6040 ;
  END
END ISOLORAOX8_LVT

MACRO ISOLORX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.216 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4910 0.5830 0.6630 0.6330 ;
        RECT 0.5530 0.5530 0.6630 0.5830 ;
        RECT 0.5530 0.6330 0.6630 0.6630 ;
    END
    ANTENNAGATEAREA 0.0306 ;
  END D

  PIN ISO
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5830 0.4210 0.6330 ;
        RECT 0.2490 0.5530 0.3590 0.5830 ;
        RECT 0.2490 0.6330 0.3590 0.6630 ;
    END
    ANTENNAGATEAREA 0.0306 ;
  END ISO

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8870 0.4730 1.0430 0.5230 ;
        RECT 0.8870 0.1270 0.9370 0.4730 ;
        RECT 0.9930 0.5230 1.0430 0.5530 ;
        RECT 0.9930 0.5530 1.1190 0.6630 ;
        RECT 0.9930 0.6630 1.0430 0.8610 ;
        RECT 0.8870 0.8610 1.0430 0.9110 ;
        RECT 0.8870 0.9110 0.9370 1.5540 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.2160 0.0300 ;
        RECT 0.4310 0.0300 0.4810 0.2090 ;
        RECT 0.7350 0.0300 0.7850 0.3010 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.2160 1.7020 ;
        RECT 0.2790 0.8150 0.3290 1.6420 ;
        RECT 0.7350 0.9170 0.7850 1.6420 ;
    END
  END VDD
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.3310 1.7730 ;
    LAYER M1 ;
      RECT 0.7420 0.6580 0.8770 0.7080 ;
      RECT 0.2790 0.3810 0.7330 0.4310 ;
      RECT 0.5830 0.7640 0.7320 0.8140 ;
      RECT 0.7130 0.3810 0.7630 0.8140 ;
      RECT 0.2790 0.1270 0.3290 0.4170 ;
      RECT 0.5830 0.1270 0.6330 0.4170 ;
      RECT 0.5830 0.7640 0.6330 1.5540 ;
    LAYER PO ;
      RECT 0.5170 0.0770 0.5470 1.6040 ;
      RECT 0.3650 0.0770 0.3950 1.6040 ;
      RECT 0.6690 0.0770 0.6990 1.6040 ;
      RECT 0.2130 0.0770 0.2430 1.6040 ;
      RECT 0.8210 0.0770 0.8510 1.6040 ;
      RECT 0.0610 0.0770 0.0910 1.6040 ;
      RECT 0.9730 0.0770 1.0030 1.6040 ;
      RECT 1.1250 0.0770 1.1550 1.6040 ;
  END
END ISOLORX1_LVT

MACRO ISOLORX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.368 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4910 0.5830 0.6630 0.6330 ;
        RECT 0.5530 0.5530 0.6630 0.5830 ;
        RECT 0.5530 0.6330 0.6630 0.6630 ;
    END
    ANTENNAGATEAREA 0.0306 ;
  END D

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8870 0.7860 1.2110 0.8360 ;
        RECT 0.8870 0.8360 0.9370 1.5560 ;
        RECT 1.1610 0.6630 1.2110 0.7860 ;
        RECT 1.1610 0.6030 1.2710 0.6630 ;
        RECT 0.8870 0.5530 1.2710 0.6030 ;
        RECT 0.8870 0.2080 0.9370 0.5530 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.3680 1.7020 ;
        RECT 1.0390 0.9220 1.0890 1.6420 ;
        RECT 0.7350 0.9220 0.7850 1.6420 ;
        RECT 0.2790 0.7380 0.3290 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.3680 0.0300 ;
        RECT 0.7350 0.0300 0.7850 0.3170 ;
        RECT 1.0390 0.0300 1.0890 0.3170 ;
        RECT 0.4310 0.0300 0.4810 0.3170 ;
    END
  END VSS

  PIN ISO
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.3590 0.5830 ;
        RECT 0.2490 0.5830 0.4210 0.6330 ;
        RECT 0.2490 0.6330 0.3590 0.6630 ;
    END
    ANTENNAGATEAREA 0.0306 ;
  END ISO
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.4830 1.7730 ;
    LAYER M1 ;
      RECT 0.7360 0.6600 1.0290 0.7100 ;
      RECT 0.2790 0.1430 0.3290 0.4330 ;
      RECT 0.5830 0.8000 0.6330 1.5560 ;
      RECT 0.5830 0.1430 0.6330 0.4330 ;
      RECT 0.5830 0.8000 0.7630 0.8500 ;
      RECT 0.2780 0.4320 0.7630 0.4820 ;
      RECT 0.7130 0.4570 0.7630 0.8500 ;
    LAYER PO ;
      RECT 1.1250 0.0930 1.1550 1.6060 ;
      RECT 0.9730 0.0930 1.0030 1.6060 ;
      RECT 0.8210 0.0930 0.8510 1.6060 ;
      RECT 1.2770 0.0930 1.3070 1.6060 ;
      RECT 0.0610 0.0930 0.0910 1.6060 ;
      RECT 0.2130 0.0930 0.2430 1.6060 ;
      RECT 0.6690 0.0930 0.6990 1.6060 ;
      RECT 0.3650 0.0930 0.3950 1.6060 ;
      RECT 0.5170 0.0930 0.5470 1.6060 ;
  END
END ISOLORX2_LVT

MACRO ISOLORX4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.672 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.6720 1.7020 ;
        RECT 0.2790 0.7360 0.3290 1.6420 ;
        RECT 1.3430 0.9200 1.3930 1.6420 ;
        RECT 0.7350 0.9200 0.7850 1.6420 ;
        RECT 1.0390 0.9200 1.0890 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.6720 0.0300 ;
        RECT 0.4310 0.0300 0.4810 0.3170 ;
        RECT 1.3430 0.0300 1.3930 0.4090 ;
        RECT 1.0390 0.0300 1.0890 0.4090 ;
        RECT 0.7350 0.0300 0.7850 0.3170 ;
    END
  END VSS

  PIN ISO
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5830 0.4210 0.6330 ;
        RECT 0.2490 0.5530 0.3590 0.5830 ;
        RECT 0.2490 0.6330 0.3590 0.6630 ;
    END
    ANTENNAGATEAREA 0.0306 ;
  END ISO

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4910 0.5830 0.6630 0.6330 ;
        RECT 0.5530 0.6330 0.6630 0.6630 ;
        RECT 0.5530 0.5530 0.6630 0.5830 ;
    END
    ANTENNAGATEAREA 0.0306 ;
  END D

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8870 0.1430 0.9370 0.5450 ;
        RECT 0.8870 0.5450 1.4680 0.5530 ;
        RECT 0.8870 0.5530 1.5750 0.5950 ;
        RECT 1.1910 0.1430 1.2410 0.5450 ;
        RECT 1.4180 0.5950 1.5750 0.6630 ;
        RECT 1.4180 0.6630 1.4680 0.7580 ;
        RECT 0.8870 0.7580 1.4680 0.8080 ;
        RECT 1.1910 0.8080 1.2410 1.5540 ;
        RECT 0.8870 0.8080 0.9370 1.5540 ;
    END
    ANTENNADIFFAREA 0.2976 ;
  END Q
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.7870 1.7730 ;
    LAYER M1 ;
      RECT 0.7500 0.6580 1.3330 0.7080 ;
      RECT 0.5830 0.8340 0.6330 1.5540 ;
      RECT 0.5830 0.1430 0.6330 0.4510 ;
      RECT 0.5830 0.7950 0.7630 0.8450 ;
      RECT 0.2780 0.4260 0.7630 0.4760 ;
      RECT 0.7130 0.4520 0.7630 0.8450 ;
      RECT 0.2790 0.1430 0.3290 0.4510 ;
    LAYER PO ;
      RECT 0.2130 0.0930 0.2430 1.6040 ;
      RECT 1.5810 0.0930 1.6110 1.6040 ;
      RECT 1.2770 0.0930 1.3070 1.6040 ;
      RECT 0.3650 0.0930 0.3950 1.6040 ;
      RECT 0.6690 0.0930 0.6990 1.6040 ;
      RECT 1.4290 0.0930 1.4590 1.6040 ;
      RECT 0.5170 0.0930 0.5470 1.6040 ;
      RECT 0.0610 0.0930 0.0910 1.6040 ;
      RECT 1.1250 0.0930 1.1550 1.6040 ;
      RECT 0.9730 0.0930 1.0030 1.6040 ;
      RECT 0.8210 0.0930 0.8510 1.6040 ;
  END
END ISOLORX4_LVT

MACRO ISOLORX8_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.584 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.5840 0.0300 ;
        RECT 0.4310 0.0300 0.4810 0.2960 ;
        RECT 1.1910 0.0300 1.2410 0.3980 ;
        RECT 1.4950 0.0300 1.5450 0.3980 ;
        RECT 2.1030 0.0300 2.1530 0.3980 ;
        RECT 1.7990 0.0300 1.8490 0.3980 ;
        RECT 0.7350 0.0300 0.7850 0.2960 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.5830 0.5730 0.6330 ;
        RECT 0.4010 0.6330 0.5110 0.6630 ;
        RECT 0.4010 0.5530 0.5110 0.5830 ;
    END
    ANTENNAGATEAREA 0.0612 ;
  END D

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3750 0.5410 2.4250 0.5530 ;
        RECT 2.3750 0.5530 2.4870 0.6630 ;
        RECT 1.0390 0.4910 2.4250 0.5410 ;
        RECT 2.3750 0.6630 2.4250 0.8450 ;
        RECT 1.9510 0.1150 2.0010 0.4910 ;
        RECT 2.2550 0.1150 2.3050 0.4910 ;
        RECT 1.0390 0.1150 1.0890 0.4910 ;
        RECT 1.3430 0.1150 1.3930 0.4910 ;
        RECT 1.6470 0.1150 1.6970 0.4910 ;
        RECT 2.3750 0.3320 2.4250 0.4910 ;
        RECT 1.0390 0.8450 2.4250 0.8950 ;
        RECT 2.2550 0.8950 2.3050 1.5440 ;
        RECT 1.0390 0.8950 1.0890 1.5440 ;
        RECT 1.9510 0.8950 2.0010 1.5440 ;
        RECT 1.3430 0.8950 1.3930 1.5440 ;
        RECT 1.6470 0.8950 1.6970 1.5440 ;
    END
    ANTENNADIFFAREA 0.6952 ;
  END Q

  PIN ISO
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6430 0.5830 0.8770 0.6330 ;
        RECT 0.7050 0.6330 0.8150 0.6630 ;
        RECT 0.7050 0.5530 0.8150 0.5830 ;
    END
    ANTENNAGATEAREA 0.0612 ;
  END ISO

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.5840 1.7020 ;
        RECT 1.7990 1.0020 1.8490 1.6420 ;
        RECT 2.1030 1.0020 2.1530 1.6420 ;
        RECT 1.4950 1.0020 1.5450 1.6420 ;
        RECT 1.1910 1.0020 1.2410 1.6420 ;
        RECT 0.7350 1.0120 0.7850 1.6420 ;
    END
  END VDD
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 2.7170 1.7730 ;
    LAYER M1 ;
      RECT 0.8870 0.8910 0.9370 1.5540 ;
      RECT 0.5830 0.8410 0.9370 0.8910 ;
      RECT 0.5830 0.8910 0.6330 1.5340 ;
      RECT 0.2790 1.5340 0.6330 1.5840 ;
      RECT 0.2790 0.8280 0.3290 1.5340 ;
      RECT 0.9310 0.5910 2.2450 0.6410 ;
      RECT 0.4310 0.7900 0.4810 1.4620 ;
      RECT 0.2790 0.1220 0.3290 0.4320 ;
      RECT 0.5830 0.1220 0.6330 0.4320 ;
      RECT 0.9310 0.4820 0.9810 0.5910 ;
      RECT 0.9310 0.6410 0.9810 0.7400 ;
      RECT 0.2790 0.4320 0.9810 0.4820 ;
      RECT 0.4310 0.7400 0.9810 0.7900 ;
      RECT 0.8870 0.1220 0.9370 0.4320 ;
    LAYER PO ;
      RECT 0.5170 0.0720 0.5470 1.6040 ;
      RECT 0.3650 0.0720 0.3950 1.6040 ;
      RECT 0.9730 0.0720 1.0030 1.6040 ;
      RECT 0.2130 0.0720 0.2430 1.6040 ;
      RECT 2.4930 0.0720 2.5230 1.6040 ;
      RECT 0.0610 0.0720 0.0910 1.6040 ;
      RECT 1.7330 0.0720 1.7630 1.6040 ;
      RECT 1.1250 0.0720 1.1550 1.6040 ;
      RECT 2.0370 0.0720 2.0670 1.6040 ;
      RECT 2.1890 0.0720 2.2190 1.6040 ;
      RECT 2.3410 0.0720 2.3710 1.6040 ;
      RECT 1.8850 0.0720 1.9150 1.6040 ;
      RECT 1.5810 0.0720 1.6110 1.6040 ;
      RECT 1.4290 0.0720 1.4590 1.6040 ;
      RECT 1.2770 0.0720 1.3070 1.6040 ;
      RECT 0.8210 0.0720 0.8510 1.6040 ;
      RECT 0.6690 0.0720 0.6990 1.6040 ;
  END
END ISOLORX8_LVT

MACRO LARX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.344 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9630 0.8570 1.1190 0.9670 ;
        RECT 0.9630 0.6830 1.0130 0.8570 ;
    END
    ANTENNAGATEAREA 0.0285 ;
  END D

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.3440 0.0300 ;
        RECT 2.8630 0.0300 2.9130 0.2200 ;
        RECT 0.4310 0.0300 0.4810 0.4500 ;
        RECT 0.5830 0.0300 0.6330 0.4500 ;
        RECT 2.5590 0.0300 2.6090 0.3180 ;
        RECT 0.8710 0.3180 2.6090 0.3680 ;
    END
  END VSS

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.7110 1.0690 3.0950 1.1190 ;
        RECT 2.9850 1.0090 3.0950 1.0690 ;
        RECT 2.7110 1.1190 2.7610 1.5460 ;
        RECT 3.0450 0.3590 3.0950 1.0090 ;
        RECT 2.7110 0.3090 3.0950 0.3590 ;
        RECT 2.7110 0.1480 2.7610 0.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.3440 1.7020 ;
        RECT 2.8630 1.1700 2.9130 1.6420 ;
        RECT 0.4910 1.3280 0.5410 1.6420 ;
        RECT 2.5990 1.3780 2.6490 1.6420 ;
        RECT 0.4310 1.2780 1.1050 1.3280 ;
        RECT 1.6310 1.3280 2.6490 1.3780 ;
        RECT 0.4310 0.7750 0.4810 1.2780 ;
        RECT 0.5830 0.7750 0.6330 1.2780 ;
    END
  END VDD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.1380 1.1610 3.2480 1.2210 ;
        RECT 3.0150 1.2210 3.2480 1.2710 ;
        RECT 3.1970 0.2040 3.2470 1.1610 ;
        RECT 3.0150 1.2710 3.0650 1.5460 ;
        RECT 2.9990 0.1540 3.2470 0.2040 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 1.4240 0.4210 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0990 0.5530 1.2710 0.6660 ;
    END
    ANTENNAGATEAREA 0.0465 ;
  END RSTB
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 3.4590 1.7730 ;
    LAYER M1 ;
      RECT 1.1750 0.4180 1.3930 0.4680 ;
      RECT 1.3430 0.4680 1.3930 1.1780 ;
      RECT 1.3430 1.2280 1.3930 1.3500 ;
      RECT 1.1910 1.0350 1.2410 1.1780 ;
      RECT 0.8870 1.1780 1.3930 1.2280 ;
      RECT 0.8870 1.0350 0.9370 1.1780 ;
      RECT 1.7830 0.5180 1.9010 0.5680 ;
      RECT 1.8510 0.5680 1.9010 0.6040 ;
      RECT 1.8510 0.6040 2.8590 0.6540 ;
      RECT 2.1430 0.6540 2.1930 0.8780 ;
      RECT 1.7830 0.8780 2.1930 0.9280 ;
      RECT 1.4950 0.4180 2.0170 0.4680 ;
      RECT 1.6680 0.4680 1.7180 0.6180 ;
      RECT 1.6680 0.6180 1.7890 0.6680 ;
      RECT 1.4950 1.1780 2.0220 1.2280 ;
      RECT 1.4950 0.4680 1.5450 1.1780 ;
      RECT 1.4950 1.2280 1.5450 1.3500 ;
      RECT 0.7350 0.0960 2.2550 0.1460 ;
      RECT 0.7350 0.5180 0.8610 0.5680 ;
      RECT 0.8110 0.5680 0.8610 0.7180 ;
      RECT 0.7350 0.7180 0.8610 0.7680 ;
      RECT 0.7350 0.1460 0.7850 0.5180 ;
      RECT 0.7350 0.7680 0.7850 0.9140 ;
      RECT 0.2790 0.6180 0.7250 0.6680 ;
      RECT 0.2790 0.6680 0.3290 1.3150 ;
      RECT 0.2790 0.1820 0.3290 0.6180 ;
      RECT 1.0990 1.4280 2.5490 1.4780 ;
      RECT 2.0870 0.4180 2.9890 0.4680 ;
      RECT 2.9390 0.4680 2.9890 0.8060 ;
      RECT 2.5750 0.8060 2.9890 0.8560 ;
      RECT 2.5750 0.8560 2.6250 1.1780 ;
      RECT 2.0870 1.1780 2.6250 1.2280 ;
      RECT 0.6380 1.5280 1.6370 1.5780 ;
      RECT 1.5550 0.1960 2.0930 0.2460 ;
      RECT 2.0100 1.5280 2.2450 1.5780 ;
    LAYER PO ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 1.2770 0.0680 1.3070 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 1.4290 0.0680 1.4590 0.6420 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 2.0370 0.0680 2.0670 0.6420 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 2.0370 1.0320 2.0670 1.6060 ;
      RECT 1.4290 1.0320 1.4590 1.6060 ;
  END
END LARX1_LVT

MACRO LARX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.648 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9630 0.8570 1.1190 0.9670 ;
        RECT 0.9630 0.6830 1.0130 0.8570 ;
    END
    ANTENNAGATEAREA 0.0285 ;
  END D

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.6480 0.0300 ;
        RECT 0.4310 0.0300 0.4810 0.4500 ;
        RECT 0.5830 0.0300 0.6330 0.4500 ;
        RECT 2.7110 0.0300 2.7610 0.2200 ;
        RECT 3.0150 0.0300 3.0650 0.2200 ;
        RECT 3.3190 0.0300 3.3690 0.2200 ;
        RECT 2.5590 0.0300 2.6090 0.3180 ;
        RECT 0.8710 0.3180 2.6090 0.3680 ;
    END
  END VSS

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8630 1.1190 2.9130 1.5460 ;
        RECT 2.8630 1.0690 3.4090 1.1190 ;
        RECT 3.2890 1.0090 3.4090 1.0690 ;
        RECT 3.3590 0.4540 3.4090 1.0090 ;
        RECT 2.8630 0.4040 3.4090 0.4540 ;
        RECT 2.8630 0.1480 2.9130 0.4040 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.6480 1.7020 ;
        RECT 2.7110 1.1700 2.7610 1.6420 ;
        RECT 3.0150 1.1700 3.0650 1.6420 ;
        RECT 3.3190 1.3720 3.3690 1.6420 ;
        RECT 0.4910 1.3280 0.5410 1.6420 ;
        RECT 2.5990 1.3780 2.6490 1.6420 ;
        RECT 0.4310 1.2780 1.1050 1.3280 ;
        RECT 1.6310 1.3280 2.6490 1.3780 ;
        RECT 0.4310 0.7750 0.4810 1.2780 ;
        RECT 0.5830 0.7750 0.6330 1.2780 ;
    END
  END VDD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.1670 1.2210 3.5860 1.2710 ;
        RECT 3.1670 1.2710 3.2170 1.5460 ;
        RECT 3.4410 1.2710 3.5860 1.4230 ;
        RECT 3.5360 0.3540 3.5860 1.2210 ;
        RECT 3.1510 0.3040 3.5860 0.3540 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 1.4240 0.4210 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0990 0.5530 1.2710 0.6660 ;
    END
    ANTENNAGATEAREA 0.0465 ;
  END RSTB
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 3.7630 1.7730 ;
    LAYER M1 ;
      RECT 1.1750 0.4180 1.3930 0.4680 ;
      RECT 1.3430 0.4680 1.3930 1.1780 ;
      RECT 1.3430 1.2280 1.3930 1.3500 ;
      RECT 1.1910 1.0350 1.2410 1.1780 ;
      RECT 0.8870 1.1780 1.3930 1.2280 ;
      RECT 0.8870 1.0350 0.9370 1.1780 ;
      RECT 1.7830 0.5180 1.9010 0.5680 ;
      RECT 1.8510 0.5680 1.9010 0.6040 ;
      RECT 1.8510 0.6040 3.0050 0.6540 ;
      RECT 2.1430 0.6540 2.1930 0.8780 ;
      RECT 1.7830 0.8780 2.1930 0.9280 ;
      RECT 1.4950 0.4180 2.0170 0.4680 ;
      RECT 1.6680 0.4680 1.7180 0.6180 ;
      RECT 1.6680 0.6180 1.7890 0.6680 ;
      RECT 1.4950 1.1780 2.0220 1.2280 ;
      RECT 1.4950 0.4680 1.5450 1.1780 ;
      RECT 1.4950 1.2280 1.5450 1.3500 ;
      RECT 0.7350 0.0960 2.2550 0.1460 ;
      RECT 0.7350 0.5180 0.8610 0.5680 ;
      RECT 0.8110 0.5680 0.8610 0.7180 ;
      RECT 0.7350 0.7180 0.8610 0.7680 ;
      RECT 0.7350 0.1460 0.7850 0.5180 ;
      RECT 0.7350 0.7680 0.7850 0.9140 ;
      RECT 3.0910 0.6040 3.3090 0.6540 ;
      RECT 3.0910 0.5540 3.1410 0.6040 ;
      RECT 3.0910 0.6540 3.1410 0.8060 ;
      RECT 2.0870 0.5040 3.1410 0.5540 ;
      RECT 2.5750 0.8060 3.1410 0.8560 ;
      RECT 2.5750 0.8560 2.6250 1.1780 ;
      RECT 2.0870 1.1780 2.6250 1.2280 ;
      RECT 0.2790 0.6180 0.7250 0.6680 ;
      RECT 0.2790 0.6680 0.3290 1.3150 ;
      RECT 0.2790 0.1820 0.3290 0.6180 ;
      RECT 1.0990 1.4280 2.5490 1.4780 ;
      RECT 0.6380 1.5280 1.6370 1.5780 ;
      RECT 1.5550 0.1960 2.0930 0.2460 ;
      RECT 2.0100 1.5280 2.2450 1.5780 ;
    LAYER PO ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 1.2770 0.0680 1.3070 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 1.4290 0.0680 1.4590 0.6420 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 2.0370 0.0680 2.0670 0.6420 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 2.0370 1.0320 2.0670 1.6060 ;
      RECT 1.4290 1.0320 1.4590 1.6060 ;
  END
END LARX2_LVT

MACRO LASRNX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.344 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9470 0.7880 1.1190 0.9670 ;
    END
    ANTENNAGATEAREA 0.0261 ;
  END D

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.3440 0.0300 ;
        RECT 0.4310 0.0300 0.4810 0.4500 ;
        RECT 0.5830 0.0300 0.6330 0.4500 ;
        RECT 2.2550 0.0300 2.3050 0.2440 ;
        RECT 3.0550 0.0300 3.1050 0.2330 ;
        RECT 0.8870 0.2440 2.7610 0.2940 ;
        RECT 3.0150 0.2330 3.1050 0.2830 ;
        RECT 0.8870 0.2940 0.9370 0.4210 ;
        RECT 2.7110 0.2940 2.7610 0.3540 ;
        RECT 3.0150 0.2830 3.0650 0.6140 ;
    END
  END VSS

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8630 0.2770 2.9130 0.7050 ;
        RECT 2.8630 0.7050 3.0950 0.7550 ;
        RECT 2.9850 0.7550 3.0950 0.8150 ;
        RECT 2.8630 0.7550 2.9130 1.5460 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.3440 1.7020 ;
        RECT 3.0150 1.1700 3.0650 1.6420 ;
        RECT 0.4910 1.3540 0.5410 1.6420 ;
        RECT 2.7510 1.3780 2.8010 1.6420 ;
        RECT 0.4310 1.3040 1.1050 1.3540 ;
        RECT 2.1280 1.3280 2.8010 1.3780 ;
        RECT 0.4310 1.0880 0.4810 1.3040 ;
        RECT 0.5830 1.1010 0.6330 1.3040 ;
        RECT 2.1280 1.2430 2.1780 1.3280 ;
        RECT 1.7830 1.1930 2.1780 1.2430 ;
    END
  END VDD

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7690 1.3130 1.9230 1.4230 ;
    END
    ANTENNAGATEAREA 0.0261 ;
  END SETB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 1.4240 0.4210 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0990 0.5530 1.2710 0.6660 ;
    END
    ANTENNAGATEAREA 0.0441 ;
  END RSTB
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 3.4590 1.7730 ;
      RECT 0.5240 0.6680 0.8410 0.6790 ;
    LAYER M1 ;
      RECT 1.9510 0.6040 2.5520 0.6540 ;
      RECT 1.9510 0.4800 2.0010 0.6040 ;
      RECT 2.2950 0.6540 2.3450 0.8780 ;
      RECT 1.6300 0.8780 2.3450 0.9280 ;
      RECT 1.4550 0.6060 1.5450 0.6560 ;
      RECT 1.4950 0.4300 1.5450 0.6060 ;
      RECT 1.4550 0.6560 1.5050 1.0010 ;
      RECT 1.4950 0.3800 2.1530 0.4300 ;
      RECT 1.4550 1.0010 2.1740 1.0510 ;
      RECT 2.1030 0.4300 2.1530 0.5540 ;
      RECT 1.7980 0.4300 1.8480 0.6180 ;
      RECT 1.7070 0.6180 1.8480 0.6680 ;
      RECT 0.7350 0.0960 2.1240 0.1460 ;
      RECT 0.7350 0.5180 0.8610 0.5680 ;
      RECT 0.8110 0.5680 0.8610 0.7180 ;
      RECT 0.7350 0.7180 0.8610 0.7680 ;
      RECT 0.7350 0.1460 0.7850 0.5180 ;
      RECT 0.7350 0.7680 0.7850 0.9140 ;
      RECT 0.2790 0.6180 0.7250 0.6680 ;
      RECT 0.2790 0.6680 0.3290 1.3540 ;
      RECT 0.2790 0.4220 0.3290 0.6180 ;
      RECT 1.5550 0.7180 2.2450 0.7680 ;
      RECT 1.1910 1.3080 1.3930 1.3580 ;
      RECT 1.1910 1.2160 1.2410 1.3080 ;
      RECT 1.3430 0.4680 1.3930 1.3080 ;
      RECT 0.8700 1.1660 1.2410 1.2160 ;
      RECT 1.1750 0.4180 1.3930 0.4680 ;
      RECT 1.0990 1.5280 2.7010 1.5780 ;
      RECT 0.6590 1.4280 1.6370 1.4780 ;
      RECT 0.6590 1.4780 0.7090 1.5820 ;
      RECT 2.2390 0.4090 2.7770 0.4590 ;
      RECT 2.7270 0.4590 2.7770 1.1180 ;
      RECT 2.2390 1.1180 2.7770 1.1680 ;
      RECT 2.0100 1.4280 2.2450 1.4780 ;
      RECT 2.4670 0.0960 3.0050 0.1460 ;
    LAYER PO ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 1.2770 0.0680 1.3070 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 2.1890 0.9320 2.2190 1.6060 ;
      RECT 1.4290 0.0680 1.4590 0.6420 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 2.1890 0.0680 2.2190 0.7960 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 1.4290 0.8820 1.4590 1.6060 ;
  END
END LASRNX1_LVT

MACRO LASRNX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.496 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9470 0.7880 1.1190 0.9670 ;
    END
    ANTENNAGATEAREA 0.0261 ;
  END D

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.4960 0.0300 ;
        RECT 0.4310 0.0300 0.4810 0.4500 ;
        RECT 0.5830 0.0300 0.6330 0.4500 ;
        RECT 3.2070 0.0300 3.2570 0.2330 ;
        RECT 2.2550 0.0300 2.3050 0.2440 ;
        RECT 3.0150 0.2330 3.2570 0.2830 ;
        RECT 0.8870 0.2440 2.7610 0.2940 ;
        RECT 3.0150 0.2830 3.0650 0.6140 ;
        RECT 0.8870 0.2940 0.9370 0.4210 ;
        RECT 2.7110 0.2940 2.7610 0.3540 ;
    END
  END VSS

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9850 0.7550 3.0950 0.8150 ;
        RECT 2.8630 0.7050 3.2170 0.7550 ;
        RECT 3.1670 0.7550 3.2170 1.5460 ;
        RECT 3.1670 0.3680 3.2170 0.7050 ;
        RECT 2.8630 0.2770 2.9130 0.7050 ;
        RECT 2.8630 0.7550 2.9130 1.5460 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.4960 1.7020 ;
        RECT 3.0150 0.9120 3.0650 1.6420 ;
        RECT 0.4910 1.3540 0.5410 1.6420 ;
        RECT 2.7510 1.3780 2.8010 1.6420 ;
        RECT 0.4310 1.3040 1.1050 1.3540 ;
        RECT 2.1280 1.3280 2.8010 1.3780 ;
        RECT 0.4310 1.0880 0.4810 1.3040 ;
        RECT 0.5830 1.1010 0.6330 1.3040 ;
        RECT 2.1280 1.2430 2.1780 1.3280 ;
        RECT 1.7830 1.1930 2.1780 1.2430 ;
    END
  END VDD

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7690 1.3130 1.9230 1.4230 ;
    END
    ANTENNAGATEAREA 0.0261 ;
  END SETB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 1.4240 0.4210 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0990 0.5530 1.2710 0.6660 ;
    END
    ANTENNAGATEAREA 0.0441 ;
  END RSTB
  OBS
    LAYER NWELL ;
      RECT 0.5320 0.6690 0.8360 0.6790 ;
      RECT -0.1150 0.6790 3.6110 1.7730 ;
    LAYER M1 ;
      RECT 1.9510 0.6040 2.5520 0.6540 ;
      RECT 1.9510 0.4800 2.0010 0.6040 ;
      RECT 2.2950 0.6540 2.3450 0.8780 ;
      RECT 1.6300 0.8780 2.3450 0.9280 ;
      RECT 1.4550 0.6060 1.5450 0.6560 ;
      RECT 1.4950 0.4300 1.5450 0.6060 ;
      RECT 1.4550 0.6560 1.5050 1.0010 ;
      RECT 1.4950 0.3800 2.1530 0.4300 ;
      RECT 1.4550 1.0010 2.1740 1.0510 ;
      RECT 2.1030 0.4300 2.1530 0.5540 ;
      RECT 1.7980 0.4300 1.8480 0.6180 ;
      RECT 1.7070 0.6180 1.8480 0.6680 ;
      RECT 0.7350 0.0960 2.1240 0.1460 ;
      RECT 0.7350 0.5180 0.8610 0.5680 ;
      RECT 0.8110 0.5680 0.8610 0.7180 ;
      RECT 0.7350 0.7180 0.8610 0.7680 ;
      RECT 0.7350 0.1460 0.7850 0.5180 ;
      RECT 0.7350 0.7680 0.7850 0.9140 ;
      RECT 0.2790 0.6180 0.7250 0.6680 ;
      RECT 0.2790 0.6680 0.3290 1.3540 ;
      RECT 0.2790 0.4220 0.3290 0.6180 ;
      RECT 2.4670 0.0960 3.1570 0.1460 ;
      RECT 1.5550 0.7180 2.2450 0.7680 ;
      RECT 1.1910 1.3080 1.3930 1.3580 ;
      RECT 1.1910 1.2160 1.2410 1.3080 ;
      RECT 1.3430 0.4680 1.3930 1.3080 ;
      RECT 0.8700 1.1660 1.2410 1.2160 ;
      RECT 1.1750 0.4180 1.3930 0.4680 ;
      RECT 1.0990 1.5280 2.7010 1.5780 ;
      RECT 0.6590 1.4280 1.6370 1.4780 ;
      RECT 0.6590 1.4780 0.7090 1.5760 ;
      RECT 2.2390 0.4090 2.7770 0.4590 ;
      RECT 2.7270 0.4590 2.7770 1.1180 ;
      RECT 2.2390 1.1180 2.7770 1.1680 ;
      RECT 2.0100 1.4280 2.2450 1.4780 ;
    LAYER PO ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 1.2770 0.0680 1.3070 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 2.1890 0.9320 2.2190 1.6060 ;
      RECT 1.4290 0.0680 1.4590 0.6420 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 2.1890 0.0680 2.2190 0.7960 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 1.4290 0.8820 1.4590 1.6060 ;
  END
END LASRNX2_LVT

MACRO LASRQX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.344 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9470 0.7880 1.1190 0.9670 ;
    END
    ANTENNAGATEAREA 0.0285 ;
  END D

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.3440 0.0300 ;
        RECT 0.4310 0.0300 0.4810 0.4500 ;
        RECT 0.5830 0.0300 0.6330 0.4500 ;
        RECT 2.8630 0.0300 2.9130 0.4880 ;
        RECT 2.2550 0.0300 2.3050 0.2440 ;
        RECT 0.8870 0.2440 2.7610 0.2940 ;
        RECT 0.8870 0.2940 0.9370 0.4210 ;
        RECT 2.7110 0.2940 2.7610 0.3540 ;
    END
  END VSS

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9850 0.7050 3.1850 0.8150 ;
        RECT 3.0150 0.8150 3.0650 1.5460 ;
        RECT 3.1350 0.5230 3.1850 0.7050 ;
        RECT 3.0150 0.4730 3.1850 0.5230 ;
        RECT 3.0150 0.2770 3.0650 0.4730 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.3440 1.7020 ;
        RECT 2.8630 1.1700 2.9130 1.6420 ;
        RECT 0.4910 1.3540 0.5410 1.6420 ;
        RECT 2.7510 1.3780 2.8010 1.6420 ;
        RECT 0.4310 1.3040 1.1050 1.3540 ;
        RECT 2.1280 1.3280 2.8010 1.3780 ;
        RECT 0.4310 1.0880 0.4810 1.3040 ;
        RECT 0.5830 1.1010 0.6330 1.3040 ;
        RECT 2.1280 1.2530 2.1780 1.3280 ;
        RECT 1.7830 1.2030 2.1780 1.2530 ;
    END
  END VDD

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7690 1.3130 1.9230 1.4540 ;
    END
    ANTENNAGATEAREA 0.0285 ;
  END SETB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 1.4240 0.4210 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0990 0.5530 1.2710 0.6660 ;
    END
    ANTENNAGATEAREA 0.0465 ;
  END RSTB
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 3.4590 1.7730 ;
      RECT 0.5250 0.6680 0.8430 0.6790 ;
    LAYER M1 ;
      RECT 1.9510 0.5660 2.5520 0.6160 ;
      RECT 1.9510 0.4440 2.0010 0.5660 ;
      RECT 2.2950 0.6160 2.3450 0.8780 ;
      RECT 1.6300 0.8780 2.3450 0.9280 ;
      RECT 1.7070 0.5660 1.8480 0.6160 ;
      RECT 1.7980 0.3940 1.8480 0.5660 ;
      RECT 1.4950 0.3440 2.1690 0.3940 ;
      RECT 2.1030 0.3940 2.1530 0.5020 ;
      RECT 1.4950 0.3940 1.5450 0.5660 ;
      RECT 1.4550 0.5660 1.5450 0.6160 ;
      RECT 1.4550 0.6160 1.5050 1.1030 ;
      RECT 1.4550 1.1030 2.1740 1.1530 ;
      RECT 0.7350 0.0960 2.1240 0.1460 ;
      RECT 0.7350 0.5180 0.8610 0.5680 ;
      RECT 0.8110 0.5680 0.8610 0.7180 ;
      RECT 0.7350 0.7180 0.8610 0.7680 ;
      RECT 0.7350 0.1460 0.7850 0.5180 ;
      RECT 0.7350 0.7680 0.7850 0.9140 ;
      RECT 0.2790 0.6180 0.7250 0.6680 ;
      RECT 0.2790 0.6680 0.3290 1.3540 ;
      RECT 0.2790 0.4220 0.3290 0.6180 ;
      RECT 1.5550 0.6660 2.2450 0.7160 ;
      RECT 1.1910 1.3080 1.3930 1.3580 ;
      RECT 1.1910 1.2160 1.2410 1.3080 ;
      RECT 1.3430 0.4680 1.3930 1.3080 ;
      RECT 0.8700 1.1660 1.2410 1.2160 ;
      RECT 1.1750 0.4180 1.3930 0.4680 ;
      RECT 1.0990 1.5280 2.7010 1.5780 ;
      RECT 0.6590 1.4280 1.6370 1.4780 ;
      RECT 0.6590 1.4780 0.7090 1.5840 ;
      RECT 2.7270 0.5840 3.0050 0.6340 ;
      RECT 2.7270 0.4590 2.7770 0.5840 ;
      RECT 2.7270 0.6340 2.7770 1.1180 ;
      RECT 2.2390 0.4090 2.7770 0.4590 ;
      RECT 2.2390 1.1180 2.7770 1.1680 ;
      RECT 2.0100 1.4280 2.2450 1.4780 ;
    LAYER PO ;
      RECT 2.1890 1.0320 2.2190 1.6060 ;
      RECT 2.1890 0.0680 2.2190 0.7440 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 1.2770 0.0680 1.3070 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 1.4290 0.0680 1.4590 0.6420 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 1.4290 0.8820 1.4590 1.6060 ;
  END
END LASRQX1_LVT

MACRO LASRQX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.496 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9470 0.7880 1.1190 0.9670 ;
    END
    ANTENNAGATEAREA 0.0285 ;
  END D

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.4960 0.0300 ;
        RECT 2.8630 0.0300 2.9130 0.4880 ;
        RECT 3.1670 0.0300 3.2170 0.3520 ;
        RECT 0.4310 0.0300 0.4810 0.4500 ;
        RECT 0.5830 0.0300 0.6330 0.4500 ;
        RECT 2.2550 0.0300 2.3050 0.2440 ;
        RECT 0.8870 0.2440 2.7610 0.2940 ;
        RECT 0.8870 0.2940 0.9370 0.4210 ;
        RECT 2.7110 0.2940 2.7610 0.3540 ;
    END
  END VSS

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9850 0.7050 3.2570 0.7550 ;
        RECT 2.9850 0.7550 3.1850 0.8150 ;
        RECT 3.2070 0.5230 3.2570 0.7050 ;
        RECT 3.0150 0.8150 3.0650 1.5460 ;
        RECT 3.0150 0.4730 3.2570 0.5230 ;
        RECT 3.0150 0.2770 3.0650 0.4730 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.4960 1.7020 ;
        RECT 3.1670 1.1700 3.2170 1.6420 ;
        RECT 2.8630 1.1700 2.9130 1.6420 ;
        RECT 0.4910 1.3540 0.5410 1.6420 ;
        RECT 2.7510 1.3780 2.8010 1.6420 ;
        RECT 0.4310 1.3040 1.1050 1.3540 ;
        RECT 2.1280 1.3280 2.8010 1.3780 ;
        RECT 0.4310 1.0880 0.4810 1.3040 ;
        RECT 0.5830 1.1010 0.6330 1.3040 ;
        RECT 2.1280 1.2530 2.1780 1.3280 ;
        RECT 1.7830 1.2030 2.1780 1.2530 ;
    END
  END VDD

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7690 1.3130 1.9230 1.4540 ;
    END
    ANTENNAGATEAREA 0.0285 ;
  END SETB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 1.4240 0.4210 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0990 0.5530 1.2710 0.6660 ;
    END
    ANTENNAGATEAREA 0.0465 ;
  END RSTB
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 3.6110 1.7730 ;
      RECT 0.5320 0.6690 0.8360 0.6790 ;
    LAYER M1 ;
      RECT 1.9510 0.5660 2.5520 0.6160 ;
      RECT 1.9510 0.4440 2.0010 0.5660 ;
      RECT 2.2950 0.6160 2.3450 0.8780 ;
      RECT 1.6300 0.8780 2.3450 0.9280 ;
      RECT 1.7070 0.5660 1.8480 0.6160 ;
      RECT 1.7980 0.3940 1.8480 0.5660 ;
      RECT 1.4950 0.3440 2.1690 0.3940 ;
      RECT 2.1030 0.3940 2.1530 0.5020 ;
      RECT 1.4950 0.3940 1.5450 0.5660 ;
      RECT 1.4550 0.5660 1.5450 0.6160 ;
      RECT 1.4550 0.6160 1.5050 1.1030 ;
      RECT 1.4550 1.1030 2.1740 1.1530 ;
      RECT 0.7350 0.0960 2.1240 0.1460 ;
      RECT 0.7350 0.5180 0.8610 0.5680 ;
      RECT 0.8110 0.5680 0.8610 0.7180 ;
      RECT 0.7350 0.7180 0.8610 0.7680 ;
      RECT 0.7350 0.1460 0.7850 0.5180 ;
      RECT 0.7350 0.7680 0.7850 0.9140 ;
      RECT 0.2790 0.6180 0.7250 0.6680 ;
      RECT 0.2790 0.6680 0.3290 1.3540 ;
      RECT 0.2790 0.4220 0.3290 0.6180 ;
      RECT 2.7270 0.5840 3.1570 0.6340 ;
      RECT 2.7270 0.4590 2.7770 0.5840 ;
      RECT 2.7270 0.6340 2.7770 1.1180 ;
      RECT 2.2390 0.4090 2.7770 0.4590 ;
      RECT 2.2390 1.1180 2.7770 1.1680 ;
      RECT 1.5550 0.6660 2.2450 0.7160 ;
      RECT 1.1910 1.3080 1.3930 1.3580 ;
      RECT 1.1910 1.2160 1.2410 1.3080 ;
      RECT 1.3430 0.4680 1.3930 1.3080 ;
      RECT 0.8700 1.1660 1.2410 1.2160 ;
      RECT 1.1750 0.4180 1.3930 0.4680 ;
      RECT 1.0990 1.5280 2.7010 1.5780 ;
      RECT 0.6590 1.4280 1.6370 1.4780 ;
      RECT 0.6590 1.4780 0.7090 1.5840 ;
      RECT 2.0100 1.4280 2.2450 1.4780 ;
    LAYER PO ;
      RECT 2.1890 1.0320 2.2190 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 2.1890 0.0680 2.2190 0.7440 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 1.2770 0.0680 1.3070 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 1.4290 0.0680 1.4590 0.6420 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 1.4290 0.8820 1.4590 1.6060 ;
  END
END LASRQX2_LVT

MACRO LASRX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.496 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9470 0.7880 1.1190 0.9670 ;
    END
    ANTENNAGATEAREA 0.0261 ;
  END D

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.4960 0.0300 ;
        RECT 0.4310 0.0300 0.4810 0.4500 ;
        RECT 0.5830 0.0300 0.6330 0.4500 ;
        RECT 3.0150 0.0300 3.0650 0.2200 ;
        RECT 2.7110 0.0300 2.7610 0.2440 ;
        RECT 0.8870 0.2440 2.7610 0.2940 ;
        RECT 0.8870 0.2940 0.9370 0.4210 ;
        RECT 2.7110 0.2940 2.7610 0.3540 ;
    END
  END VSS

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8630 1.0690 3.2470 1.1190 ;
        RECT 3.1370 1.0090 3.2470 1.0690 ;
        RECT 2.8630 1.1190 2.9130 1.5460 ;
        RECT 3.1970 0.3590 3.2470 1.0090 ;
        RECT 2.8630 0.3090 3.2470 0.3590 ;
        RECT 2.8630 0.1480 2.9130 0.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.4960 1.7020 ;
        RECT 3.0150 1.1700 3.0650 1.6420 ;
        RECT 0.4910 1.3540 0.5410 1.6420 ;
        RECT 2.7510 1.3780 2.8010 1.6420 ;
        RECT 0.4310 1.3040 1.1050 1.3540 ;
        RECT 2.1280 1.3280 2.8010 1.3780 ;
        RECT 0.4310 1.0880 0.4810 1.3040 ;
        RECT 0.5830 1.1010 0.6330 1.3040 ;
        RECT 2.1280 1.2430 2.1780 1.3280 ;
        RECT 1.7830 1.1930 2.1780 1.2430 ;
    END
  END VDD

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7690 1.3130 1.9230 1.4230 ;
    END
    ANTENNAGATEAREA 0.0261 ;
  END SETB

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2900 1.1610 3.4000 1.2210 ;
        RECT 3.1670 1.2210 3.4000 1.2710 ;
        RECT 3.3490 0.2040 3.3990 1.1610 ;
        RECT 3.1670 1.2710 3.2170 1.5460 ;
        RECT 3.1510 0.1540 3.3990 0.2040 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 1.4240 0.4210 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0990 0.5530 1.2710 0.6660 ;
    END
    ANTENNAGATEAREA 0.0441 ;
  END RSTB
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 3.6110 1.7730 ;
      RECT 0.5240 0.6680 0.8450 0.6790 ;
    LAYER M1 ;
      RECT 1.4550 0.6060 1.5450 0.6560 ;
      RECT 1.4950 0.4300 1.5450 0.6060 ;
      RECT 1.4550 0.6560 1.5050 1.0010 ;
      RECT 1.4950 0.3800 2.1530 0.4300 ;
      RECT 1.4550 1.0010 2.1740 1.0510 ;
      RECT 2.1030 0.4300 2.1530 0.5540 ;
      RECT 1.7980 0.4300 1.8480 0.6180 ;
      RECT 1.7070 0.6180 1.8480 0.6680 ;
      RECT 1.9510 0.6040 3.0110 0.6540 ;
      RECT 1.9510 0.4800 2.0010 0.6040 ;
      RECT 2.2950 0.6540 2.3450 0.8780 ;
      RECT 1.6300 0.8780 2.3450 0.9280 ;
      RECT 0.7350 0.0960 2.1240 0.1460 ;
      RECT 0.7350 0.5180 0.8610 0.5680 ;
      RECT 0.8110 0.5680 0.8610 0.7180 ;
      RECT 0.7350 0.7180 0.8610 0.7680 ;
      RECT 0.7350 0.1460 0.7850 0.5180 ;
      RECT 0.7350 0.7680 0.7850 0.9140 ;
      RECT 0.2790 0.6180 0.7250 0.6680 ;
      RECT 0.2790 0.6680 0.3290 1.3540 ;
      RECT 0.2790 0.4220 0.3290 0.6180 ;
      RECT 1.5550 0.7180 2.2450 0.7680 ;
      RECT 1.1910 1.3080 1.3930 1.3580 ;
      RECT 1.1910 1.2160 1.2410 1.3080 ;
      RECT 1.3430 0.4680 1.3930 1.3080 ;
      RECT 0.8700 1.1660 1.2410 1.2160 ;
      RECT 1.1750 0.4180 1.3930 0.4680 ;
      RECT 1.0990 1.5280 2.7010 1.5780 ;
      RECT 2.2390 0.4090 3.1410 0.4590 ;
      RECT 3.0910 0.4590 3.1410 0.8060 ;
      RECT 2.7270 0.8060 3.1410 0.8560 ;
      RECT 2.7270 0.8560 2.7770 1.1180 ;
      RECT 2.2390 1.1180 2.7770 1.1680 ;
      RECT 0.6590 1.4280 1.6370 1.4780 ;
      RECT 0.6590 1.4780 0.7090 1.5840 ;
      RECT 2.0100 1.4280 2.2450 1.4780 ;
    LAYER PO ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 1.2770 0.0680 1.3070 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 2.1890 0.9320 2.2190 1.6060 ;
      RECT 1.4290 0.0680 1.4590 0.6420 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 2.1890 0.0680 2.2190 0.7960 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 1.4290 0.8820 1.4590 1.6060 ;
  END
END LASRX1_LVT

MACRO INVX32_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.472 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6600 5.1480 0.7100 ;
        RECT 0.2490 0.7100 0.3620 0.8150 ;
    END
    ANTENNAGATEAREA 1.1712 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 5.4720 1.7020 ;
        RECT 4.9910 0.9920 5.0410 1.6420 ;
        RECT 4.6870 0.9920 4.7370 1.6420 ;
        RECT 4.3830 0.9920 4.4330 1.6420 ;
        RECT 4.0790 0.9920 4.1290 1.6420 ;
        RECT 3.7750 0.9920 3.8250 1.6420 ;
        RECT 3.4710 0.9920 3.5210 1.6420 ;
        RECT 3.1670 0.9920 3.2170 1.6420 ;
        RECT 2.8630 0.9920 2.9130 1.6420 ;
        RECT 2.5590 0.9920 2.6090 1.6420 ;
        RECT 2.2550 0.9920 2.3050 1.6420 ;
        RECT 1.9510 0.9920 2.0010 1.6420 ;
        RECT 1.6470 0.9920 1.6970 1.6420 ;
        RECT 1.0390 0.9920 1.0890 1.6420 ;
        RECT 1.3430 0.9920 1.3930 1.6420 ;
        RECT 0.7350 0.9920 0.7850 1.6420 ;
        RECT 0.4310 0.9920 0.4810 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 5.4720 0.0300 ;
        RECT 0.4310 0.0300 0.4810 0.4100 ;
        RECT 4.9910 0.0300 5.0410 0.4100 ;
        RECT 4.6870 0.0300 4.7370 0.4100 ;
        RECT 4.3830 0.0300 4.4330 0.4100 ;
        RECT 4.0790 0.0300 4.1290 0.4100 ;
        RECT 3.7750 0.0300 3.8250 0.4100 ;
        RECT 3.4710 0.0300 3.5210 0.4100 ;
        RECT 3.1670 0.0300 3.2170 0.4100 ;
        RECT 2.8630 0.0300 2.9130 0.4100 ;
        RECT 2.5590 0.0300 2.6090 0.4100 ;
        RECT 2.2550 0.0300 2.3050 0.4100 ;
        RECT 1.9510 0.0300 2.0010 0.4100 ;
        RECT 1.6470 0.0300 1.6970 0.4100 ;
        RECT 1.0390 0.0300 1.0890 0.4100 ;
        RECT 1.3430 0.0300 1.3930 0.4100 ;
        RECT 0.7350 0.0300 0.7850 0.4100 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.0150 0.9420 3.0650 1.5640 ;
        RECT 3.3190 0.9420 3.3690 1.5640 ;
        RECT 3.6230 0.9420 3.6730 1.5640 ;
        RECT 3.9270 0.9420 3.9770 1.5640 ;
        RECT 4.2310 0.9420 4.2810 1.5640 ;
        RECT 4.5350 0.9420 4.5850 1.5640 ;
        RECT 4.8390 0.9420 4.8890 1.5640 ;
        RECT 5.1430 0.9420 5.1930 1.5640 ;
        RECT 1.4950 0.9420 1.5450 1.5650 ;
        RECT 0.8870 0.9420 0.9370 1.5640 ;
        RECT 0.5830 0.9420 0.6330 1.5640 ;
        RECT 0.2790 0.9420 0.3290 1.5640 ;
        RECT 1.7990 0.9420 1.8490 1.5640 ;
        RECT 1.1910 0.9420 1.2410 1.5640 ;
        RECT 2.1030 0.9420 2.1530 1.5640 ;
        RECT 2.4070 0.9420 2.4570 1.5640 ;
        RECT 2.7110 0.9420 2.7610 1.5640 ;
        RECT 0.2790 0.8920 5.2520 0.9420 ;
        RECT 5.2020 0.6630 5.2520 0.8920 ;
        RECT 0.2790 0.5370 5.3750 0.5870 ;
        RECT 0.5830 0.1160 0.6330 0.5370 ;
        RECT 0.2790 0.1160 0.3290 0.5370 ;
        RECT 0.8870 0.1160 0.9370 0.5370 ;
        RECT 2.1030 0.1160 2.1530 0.5370 ;
        RECT 1.7990 0.1160 1.8490 0.5370 ;
        RECT 1.4950 0.1170 1.5450 0.5370 ;
        RECT 1.1910 0.1160 1.2410 0.5370 ;
        RECT 2.4070 0.1160 2.4570 0.5370 ;
        RECT 2.7110 0.1160 2.7610 0.5370 ;
        RECT 5.2020 0.5870 5.3750 0.6630 ;
        RECT 3.0150 0.1160 3.0650 0.5370 ;
        RECT 3.3190 0.1160 3.3690 0.5370 ;
        RECT 3.6230 0.1160 3.6730 0.5370 ;
        RECT 3.9270 0.1160 3.9770 0.5370 ;
        RECT 4.2310 0.1160 4.2810 0.5370 ;
        RECT 4.5350 0.1160 4.5850 0.5370 ;
        RECT 4.8390 0.1160 4.8890 0.5370 ;
        RECT 5.1430 0.1160 5.1930 0.5370 ;
    END
    ANTENNADIFFAREA 2.4808 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 5.5870 1.7730 ;
    LAYER PO ;
      RECT 5.3810 0.0690 5.4110 1.6060 ;
      RECT 5.2290 0.0690 5.2590 1.6060 ;
      RECT 5.0770 0.0690 5.1070 1.6060 ;
      RECT 4.9250 0.0690 4.9550 1.6060 ;
      RECT 4.6210 0.0690 4.6510 1.6060 ;
      RECT 4.7730 0.0690 4.8030 1.6060 ;
      RECT 4.3170 0.0690 4.3470 1.6060 ;
      RECT 4.4690 0.0690 4.4990 1.6060 ;
      RECT 4.1650 0.0690 4.1950 1.6060 ;
      RECT 4.0130 0.0690 4.0430 1.6060 ;
      RECT 3.8610 0.0690 3.8910 1.6060 ;
      RECT 3.7090 0.0690 3.7390 1.6060 ;
      RECT 3.4050 0.0690 3.4350 1.6060 ;
      RECT 3.5570 0.0690 3.5870 1.6060 ;
      RECT 2.7970 0.0690 2.8270 1.6060 ;
      RECT 2.9490 0.0690 2.9790 1.6060 ;
      RECT 2.6450 0.0690 2.6750 1.6060 ;
      RECT 3.1010 0.0690 3.1310 1.6060 ;
      RECT 3.2530 0.0690 3.2830 1.6060 ;
      RECT 1.4290 0.0690 1.4590 1.6060 ;
      RECT 1.5810 0.0690 1.6110 1.6060 ;
      RECT 1.7330 0.0690 1.7630 1.6060 ;
      RECT 2.3410 0.0690 2.3710 1.6060 ;
      RECT 2.1890 0.0690 2.2190 1.6060 ;
      RECT 2.0370 0.0690 2.0670 1.6060 ;
      RECT 1.8850 0.0690 1.9150 1.6060 ;
      RECT 2.4930 0.0690 2.5230 1.6060 ;
      RECT 1.2770 0.0690 1.3070 1.6060 ;
      RECT 1.1250 0.0690 1.1550 1.6060 ;
      RECT 0.9730 0.0690 1.0030 1.6060 ;
      RECT 0.2130 0.0690 0.2430 1.6060 ;
      RECT 0.3650 0.0690 0.3950 1.6060 ;
      RECT 0.8210 0.0690 0.8510 1.6060 ;
      RECT 0.6690 0.0690 0.6990 1.6060 ;
      RECT 0.5170 0.0690 0.5470 1.6060 ;
      RECT 0.0610 0.0690 0.0910 1.6060 ;
  END
END INVX32_LVT

MACRO INVX4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.216 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6600 0.8920 0.7100 ;
        RECT 0.2490 0.7100 0.3620 0.8150 ;
    END
    ANTENNAGATEAREA 0.1464 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.2160 1.7020 ;
        RECT 0.7350 0.9920 0.7850 1.6420 ;
        RECT 0.4310 0.9920 0.4810 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.2160 0.0300 ;
        RECT 0.7350 0.0300 0.7850 0.4100 ;
        RECT 0.4310 0.0300 0.4810 0.4100 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2790 0.5370 1.1190 0.5870 ;
        RECT 0.9420 0.5870 1.1190 0.6630 ;
        RECT 0.8870 0.1160 0.9370 0.5370 ;
        RECT 0.2790 0.1160 0.3290 0.5370 ;
        RECT 0.5830 0.1160 0.6330 0.5370 ;
        RECT 0.9420 0.6630 0.9920 0.8920 ;
        RECT 0.2790 0.8920 0.9920 0.9420 ;
        RECT 0.2790 0.9420 0.3290 1.5640 ;
        RECT 0.5830 0.9420 0.6330 1.5640 ;
        RECT 0.8870 0.9420 0.9370 1.5640 ;
    END
    ANTENNADIFFAREA 0.3976 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1120 0.6790 1.3310 1.7730 ;
    LAYER PO ;
      RECT 1.1250 0.0650 1.1550 1.6000 ;
      RECT 0.9730 0.0650 1.0030 1.6000 ;
      RECT 0.2130 0.0710 0.2430 1.6060 ;
      RECT 0.3650 0.0690 0.3950 1.6060 ;
      RECT 0.8210 0.0690 0.8510 1.6060 ;
      RECT 0.6690 0.0690 0.6990 1.6060 ;
      RECT 0.5170 0.0690 0.5470 1.6060 ;
      RECT 0.0610 0.0710 0.0910 1.6060 ;
  END
END INVX4_LVT

MACRO INVX8_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.824 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6600 1.5000 0.7100 ;
        RECT 0.2490 0.7100 0.3620 0.8150 ;
    END
    ANTENNAGATEAREA 0.2928 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.8240 1.7020 ;
        RECT 1.0390 0.9920 1.0890 1.6420 ;
        RECT 1.3430 0.9920 1.3930 1.6420 ;
        RECT 0.7350 0.9920 0.7850 1.6420 ;
        RECT 0.4310 0.9920 0.4810 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.8240 0.0300 ;
        RECT 1.0390 0.0300 1.0890 0.4100 ;
        RECT 1.3430 0.0300 1.3930 0.4100 ;
        RECT 0.7350 0.0300 0.7850 0.4100 ;
        RECT 0.4310 0.0300 0.4810 0.4100 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2790 0.5370 1.7270 0.5870 ;
        RECT 1.5510 0.5870 1.7270 0.6630 ;
        RECT 1.1910 0.1160 1.2410 0.5370 ;
        RECT 1.4950 0.1170 1.5450 0.5370 ;
        RECT 0.8870 0.1160 0.9370 0.5370 ;
        RECT 0.2790 0.1160 0.3290 0.5370 ;
        RECT 0.5830 0.1160 0.6330 0.5370 ;
        RECT 1.5510 0.6630 1.6010 0.8920 ;
        RECT 0.2790 0.8920 1.6010 0.9420 ;
        RECT 1.1910 0.9420 1.2410 1.5640 ;
        RECT 1.4950 0.9420 1.5450 1.5650 ;
        RECT 0.2790 0.9420 0.3290 1.5640 ;
        RECT 0.5830 0.9420 0.6330 1.5640 ;
        RECT 0.8870 0.9420 0.9370 1.5640 ;
    END
    ANTENNADIFFAREA 0.6952 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.9390 1.7730 ;
    LAYER PO ;
      RECT 1.4290 0.0690 1.4590 1.6060 ;
      RECT 1.5810 0.0690 1.6110 1.6060 ;
      RECT 1.7330 0.0690 1.7630 1.6060 ;
      RECT 1.2770 0.0690 1.3070 1.6060 ;
      RECT 1.1250 0.0690 1.1550 1.6060 ;
      RECT 0.9730 0.0690 1.0030 1.6060 ;
      RECT 0.2130 0.0690 0.2430 1.6060 ;
      RECT 0.3650 0.0690 0.3950 1.6060 ;
      RECT 0.8210 0.0690 0.8510 1.6060 ;
      RECT 0.6690 0.0690 0.6990 1.6060 ;
      RECT 0.5170 0.0690 0.5470 1.6060 ;
      RECT 0.0610 0.0690 0.0910 1.6060 ;
  END
END INVX8_LVT

MACRO ISOLANDAOX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.344 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.5550 1.3430 1.7890 1.3930 ;
        RECT 1.6170 1.3930 1.7270 1.4230 ;
        RECT 1.6170 1.3130 1.7270 1.3430 ;
    END
    ANTENNAGATEAREA 0.0234 ;
  END D

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.3440 1.7020 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.3440 0.0300 ;
        RECT 1.3430 0.0300 1.3930 0.3000 ;
        RECT 1.0390 0.0300 1.0890 0.3260 ;
        RECT 2.2950 0.0300 2.3450 0.2150 ;
        RECT 2.1030 0.2150 2.3450 0.2650 ;
        RECT 2.1030 0.2650 2.1530 0.3980 ;
    END
  END VSS

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 2.3770 0.7050 2.4870 0.8150 ;
        RECT 2.4070 0.6830 2.4570 0.7050 ;
        RECT 2.4070 0.8150 2.4570 0.9860 ;
        RECT 2.1030 0.9860 2.4570 1.0360 ;
        RECT 2.1030 0.6170 2.1530 0.9860 ;
        RECT 2.4070 1.0360 2.4570 1.2000 ;
        RECT 1.0370 1.2000 2.4570 1.2500 ;
        RECT 1.0390 0.6710 1.0890 1.2000 ;
        RECT 1.3430 0.8540 1.3930 1.2000 ;
        RECT 1.6470 0.8540 1.6970 1.2000 ;
    END
  END VDDG

  PIN ISO
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9470 0.4060 1.1190 0.4560 ;
        RECT 1.0090 0.3760 1.1190 0.4060 ;
        RECT 1.0090 0.4560 1.1190 0.5110 ;
    END
    ANTENNAGATEAREA 0.0186 ;
  END ISO

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9510 0.2240 2.0010 0.4600 ;
        RECT 1.9510 0.4600 2.3350 0.5100 ;
        RECT 2.2250 0.5100 2.3350 0.5110 ;
        RECT 2.2250 0.4010 2.3350 0.4600 ;
        RECT 1.9510 0.5100 2.0010 0.9760 ;
        RECT 2.2550 0.5110 2.3050 0.9360 ;
        RECT 2.2550 0.3160 2.3050 0.4010 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q
  OBS
    LAYER NWELL ;
      RECT 0.8060 0.4530 2.7110 1.0830 ;
      RECT -0.0910 1.5430 3.4590 1.7730 ;
      RECT -0.0910 0.6790 0.3460 1.5430 ;
      RECT 3.1710 0.6790 3.4590 1.5430 ;
    LAYER M1 ;
      RECT 1.4950 0.0880 1.8490 0.1380 ;
      RECT 1.7990 0.1380 1.8490 0.3000 ;
      RECT 1.4950 0.1380 1.5450 0.3500 ;
      RECT 1.1910 0.3500 1.5450 0.4000 ;
      RECT 1.1910 0.1260 1.2410 0.3500 ;
      RECT 1.7990 1.0860 2.2590 1.1360 ;
      RECT 1.1910 0.7670 1.2410 1.0180 ;
      RECT 1.4950 0.7670 1.5450 1.0280 ;
      RECT 1.7990 0.7670 1.8490 1.0860 ;
      RECT 1.1910 0.7170 1.8490 0.7670 ;
      RECT 1.6470 0.1980 1.6970 0.7170 ;
      RECT 0.8870 1.3280 1.4850 1.3780 ;
      RECT 0.8870 0.5710 0.9370 1.3280 ;
      RECT 0.8470 0.5210 0.9370 0.5710 ;
      RECT 0.8470 0.2890 0.9370 0.3390 ;
      RECT 0.8870 0.1210 0.9370 0.2890 ;
      RECT 0.8470 0.3390 0.8970 0.5210 ;
    LAYER PO ;
      RECT 1.5810 0.0710 1.6110 1.6030 ;
      RECT 1.7330 0.0710 1.7630 1.6040 ;
      RECT 2.6450 0.0720 2.6750 1.6040 ;
      RECT 0.9730 0.0710 1.0030 1.6030 ;
      RECT 1.1250 0.0710 1.1550 1.6030 ;
      RECT 0.8210 0.0710 0.8510 1.6030 ;
      RECT 2.1890 0.0720 2.2190 1.6100 ;
      RECT 0.6690 0.0710 0.6990 1.6040 ;
      RECT 2.9490 0.0720 2.9790 1.6100 ;
      RECT 0.5170 0.0710 0.5470 1.6030 ;
      RECT 2.7970 0.0720 2.8270 1.6030 ;
      RECT 1.2770 0.0710 1.3070 1.6030 ;
      RECT 1.8850 0.0720 1.9150 1.6040 ;
      RECT 2.3410 0.0710 2.3710 1.6030 ;
      RECT 1.4290 0.0710 1.4590 1.6040 ;
      RECT 2.0370 0.0720 2.0670 1.6030 ;
      RECT 2.4930 0.0720 2.5230 1.6040 ;
  END
END ISOLANDAOX1_LVT

MACRO ISOLANDAOX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.496 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7990 0.4610 2.4870 0.5110 ;
        RECT 2.4070 0.5110 2.4570 1.0280 ;
        RECT 1.7990 0.1870 1.8490 0.4610 ;
        RECT 2.3770 0.4010 2.4870 0.4610 ;
        RECT 1.7990 0.5110 1.8490 1.0280 ;
        RECT 2.1030 0.5110 2.1530 1.0280 ;
        RECT 2.1030 0.1900 2.1530 0.4610 ;
        RECT 2.4070 0.1900 2.4570 0.4010 ;
    END
    ANTENNADIFFAREA 0.1988 ;
  END Q

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 2.5290 0.7050 2.6390 0.8150 ;
        RECT 2.5590 0.6830 2.6090 0.7050 ;
        RECT 2.5590 0.8150 2.6090 1.0780 ;
        RECT 1.9510 1.0780 2.6090 1.1280 ;
        RECT 1.9510 0.6700 2.0010 1.0780 ;
        RECT 2.2550 0.6700 2.3050 1.0780 ;
        RECT 2.5590 1.1280 2.6090 1.2920 ;
        RECT 0.8850 1.2920 2.6090 1.3420 ;
        RECT 1.1910 0.8540 1.2410 1.2920 ;
        RECT 0.8870 0.6710 0.9370 1.2920 ;
        RECT 1.4950 0.8540 1.5450 1.2920 ;
    END
  END VDDG

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4030 1.4570 1.6370 1.5070 ;
        RECT 1.4650 1.5070 1.5750 1.5750 ;
    END
    ANTENNAGATEAREA 0.0234 ;
  END D

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.4960 1.7020 ;
    END
  END VDD

  PIN ISO
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7950 0.4060 0.9670 0.4560 ;
        RECT 0.8570 0.3760 0.9670 0.4060 ;
        RECT 0.8570 0.4560 0.9670 0.5110 ;
    END
    ANTENNAGATEAREA 0.0198 ;
  END ISO

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.4960 0.0300 ;
        RECT 1.1910 0.0300 1.2410 0.3260 ;
        RECT 0.8870 0.0300 0.9370 0.3260 ;
        RECT 2.4480 0.0300 2.4980 0.0880 ;
        RECT 1.9510 0.0880 2.4980 0.1380 ;
        RECT 1.9510 0.1380 2.0010 0.3720 ;
        RECT 2.2550 0.1380 2.3050 0.3720 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.0910 1.5430 3.6110 1.7730 ;
      RECT -0.0910 0.6790 0.1940 1.5430 ;
      RECT 3.3230 0.6790 3.6110 1.5430 ;
      RECT 0.6540 0.4530 2.8630 1.0830 ;
    LAYER M1 ;
      RECT 1.0390 0.3870 1.3930 0.4370 ;
      RECT 1.3430 0.1410 1.3930 0.3870 ;
      RECT 1.3430 0.0910 1.6970 0.1410 ;
      RECT 1.6470 0.1410 1.6970 0.3370 ;
      RECT 1.0390 0.1630 1.0890 0.3870 ;
      RECT 0.7350 1.3920 1.3330 1.4420 ;
      RECT 0.7350 0.5710 0.7850 1.3920 ;
      RECT 0.6950 0.5210 0.7850 0.5710 ;
      RECT 0.6950 0.2890 0.7850 0.3390 ;
      RECT 0.7350 0.1210 0.7850 0.2890 ;
      RECT 0.6950 0.3390 0.7450 0.5210 ;
      RECT 1.6470 1.1920 2.3970 1.2420 ;
      RECT 1.0390 0.7670 1.0890 1.0180 ;
      RECT 1.3430 0.7670 1.3930 1.0280 ;
      RECT 1.6470 0.7670 1.6970 1.1920 ;
      RECT 1.0390 0.7170 1.6970 0.7670 ;
      RECT 1.4950 0.1910 1.5450 0.7170 ;
    LAYER PO ;
      RECT 3.4050 0.0720 3.4350 1.6040 ;
      RECT 2.3410 0.0720 2.3710 1.6040 ;
      RECT 3.1010 0.0720 3.1310 1.6040 ;
      RECT 1.4290 0.0710 1.4590 1.6040 ;
      RECT 1.8850 0.0720 1.9150 1.6030 ;
      RECT 1.2770 0.0710 1.3070 1.6040 ;
      RECT 2.1890 0.0710 2.2190 1.6030 ;
      RECT 1.7330 0.0720 1.7630 1.6040 ;
      RECT 1.1250 0.0710 1.1550 1.6030 ;
      RECT 2.6450 0.0720 2.6750 1.6030 ;
      RECT 0.3650 0.0710 0.3950 1.6030 ;
      RECT 2.7970 0.0720 2.8270 1.6100 ;
      RECT 0.5170 0.0710 0.5470 1.6040 ;
      RECT 2.9490 0.0710 2.9790 1.6030 ;
      RECT 2.0370 0.0720 2.0670 1.6100 ;
      RECT 0.6690 0.0710 0.6990 1.6030 ;
      RECT 0.9730 0.0710 1.0030 1.6030 ;
      RECT 0.8210 0.0710 0.8510 1.6030 ;
      RECT 2.4930 0.0720 2.5230 1.6040 ;
      RECT 3.2530 0.0720 3.2830 1.6040 ;
      RECT 1.5810 0.0710 1.6110 1.6040 ;
  END
END ISOLANDAOX2_LVT

MACRO ISOLANDAOX4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.104 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 3.1370 0.7050 3.2470 0.8150 ;
        RECT 3.1670 0.6830 3.2170 0.7050 ;
        RECT 3.1670 0.8150 3.2170 1.0780 ;
        RECT 1.9510 1.0780 3.2170 1.1280 ;
        RECT 1.9510 0.6700 2.0010 1.0780 ;
        RECT 2.5590 0.6700 2.6090 1.0780 ;
        RECT 2.2550 0.6700 2.3050 1.0780 ;
        RECT 2.8630 0.6700 2.9130 1.0780 ;
        RECT 3.1670 1.1280 3.2170 1.3140 ;
        RECT 0.8850 1.3140 3.2170 1.3640 ;
        RECT 1.4950 0.8540 1.5450 1.3140 ;
        RECT 1.1910 0.8540 1.2410 1.3140 ;
        RECT 0.8870 0.6710 0.9370 1.3140 ;
    END
  END VDDG

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7990 0.4610 3.0950 0.5110 ;
        RECT 1.7990 0.2240 1.8490 0.4610 ;
        RECT 2.9850 0.4010 3.0950 0.4610 ;
        RECT 3.0150 0.5110 3.0650 1.0180 ;
        RECT 1.7990 0.5110 1.8490 1.0280 ;
        RECT 2.4070 0.5110 2.4570 1.0180 ;
        RECT 2.4070 0.2240 2.4570 0.4610 ;
        RECT 2.7110 0.5110 2.7610 1.0180 ;
        RECT 2.7110 0.2240 2.7610 0.4610 ;
        RECT 2.1030 0.5110 2.1530 1.0180 ;
        RECT 2.1030 0.2240 2.1530 0.4610 ;
        RECT 3.0150 0.2240 3.0650 0.4010 ;
    END
    ANTENNADIFFAREA 0.3476 ;
  END Q

  PIN ISO
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7950 0.4060 0.9670 0.4560 ;
        RECT 0.8570 0.4560 0.9670 0.4860 ;
        RECT 0.8570 0.3760 0.9670 0.4060 ;
    END
    ANTENNAGATEAREA 0.0186 ;
  END ISO

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.1040 0.0300 ;
        RECT 1.9510 0.0300 2.0010 0.3980 ;
        RECT 2.5590 0.0300 2.6090 0.3980 ;
        RECT 2.8630 0.0300 2.9130 0.3980 ;
        RECT 2.2550 0.0300 2.3050 0.3980 ;
        RECT 1.1910 0.0300 1.2410 0.3000 ;
        RECT 0.8870 0.0300 0.9370 0.3260 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.1040 1.7020 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4030 1.4440 1.6370 1.4940 ;
        RECT 1.4650 1.4940 1.5750 1.5750 ;
    END
    ANTENNAGATEAREA 0.0234 ;
  END D
  OBS
    LAYER NWELL ;
      RECT -0.0910 1.5430 4.2250 1.7730 ;
      RECT -0.0910 0.6790 0.1940 1.5430 ;
      RECT 3.9310 0.6790 4.2250 1.5430 ;
      RECT 0.6540 0.4530 3.4710 1.0830 ;
    LAYER M1 ;
      RECT 1.3430 0.0880 1.6970 0.1380 ;
      RECT 1.6470 0.1380 1.6970 0.3000 ;
      RECT 1.3430 0.1380 1.3930 0.3500 ;
      RECT 1.0390 0.3500 1.3930 0.4000 ;
      RECT 1.0390 0.1260 1.0890 0.3500 ;
      RECT 1.6470 1.2040 3.0050 1.2540 ;
      RECT 1.0390 0.7670 1.0890 1.0180 ;
      RECT 1.3430 0.7670 1.3930 1.0280 ;
      RECT 1.6470 0.7670 1.6970 1.2040 ;
      RECT 1.0390 0.7170 1.6970 0.7670 ;
      RECT 1.4950 0.2130 1.5450 0.7170 ;
      RECT 0.7350 1.4290 1.3330 1.4790 ;
      RECT 0.7350 0.5710 0.7850 1.4290 ;
      RECT 0.6950 0.5210 0.7850 0.5710 ;
      RECT 0.6950 0.2890 0.7850 0.3390 ;
      RECT 0.7350 0.1210 0.7850 0.2890 ;
      RECT 0.6950 0.3390 0.7450 0.5210 ;
    LAYER PO ;
      RECT 3.1010 0.0720 3.1310 1.6040 ;
      RECT 3.2530 0.0720 3.2830 1.6030 ;
      RECT 3.4050 0.0720 3.4350 1.6100 ;
      RECT 3.5570 0.0720 3.5870 1.6100 ;
      RECT 2.9490 0.0720 2.9790 1.6100 ;
      RECT 2.3410 0.0720 2.3710 1.6040 ;
      RECT 1.8850 0.0720 1.9150 1.6030 ;
      RECT 1.2770 0.0710 1.3070 1.6040 ;
      RECT 2.1890 0.0710 2.2190 1.6030 ;
      RECT 1.7330 0.0720 1.7630 1.6040 ;
      RECT 1.1250 0.0710 1.1550 1.6030 ;
      RECT 2.6450 0.0720 2.6750 1.6030 ;
      RECT 0.3650 0.0710 0.3950 1.6030 ;
      RECT 2.7970 0.0720 2.8270 1.6100 ;
      RECT 0.5170 0.0710 0.5470 1.6040 ;
      RECT 2.0370 0.0720 2.0670 1.6100 ;
      RECT 0.6690 0.0710 0.6990 1.6030 ;
      RECT 0.9730 0.0710 1.0030 1.6030 ;
      RECT 0.8210 0.0710 0.8510 1.6030 ;
      RECT 2.4930 0.0720 2.5230 1.6040 ;
      RECT 1.5810 0.0710 1.6110 1.6040 ;
      RECT 1.4290 0.0710 1.4590 1.6030 ;
  END
END ISOLANDAOX4_LVT

MACRO ISOLANDAOX8_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.32 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7990 0.4610 4.3100 0.5110 ;
        RECT 1.7990 0.1260 1.8490 0.4610 ;
        RECT 4.2000 0.4010 4.3100 0.4610 ;
        RECT 4.2310 0.5110 4.2810 1.0280 ;
        RECT 2.1030 0.5110 2.1530 1.0280 ;
        RECT 2.1030 0.1260 2.1530 0.4610 ;
        RECT 1.7990 0.5110 1.8490 1.0280 ;
        RECT 2.4070 0.5110 2.4570 1.0280 ;
        RECT 2.4070 0.1260 2.4570 0.4610 ;
        RECT 2.7110 0.5110 2.7610 1.0280 ;
        RECT 2.7110 0.1260 2.7610 0.4610 ;
        RECT 3.0150 0.5110 3.0650 1.0280 ;
        RECT 3.0150 0.1260 3.0650 0.4610 ;
        RECT 3.6230 0.5110 3.6730 1.0280 ;
        RECT 3.6230 0.1260 3.6730 0.4610 ;
        RECT 3.3190 0.5110 3.3690 1.0280 ;
        RECT 3.3190 0.1260 3.3690 0.4610 ;
        RECT 3.9270 0.5110 3.9770 1.0280 ;
        RECT 3.9270 0.1260 3.9770 0.4610 ;
        RECT 4.2310 0.1260 4.2810 0.4010 ;
    END
    ANTENNADIFFAREA 0.6452 ;
  END Q

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 4.3530 0.7050 4.4630 0.8150 ;
        RECT 4.3830 0.6830 4.4330 0.7050 ;
        RECT 4.3830 0.8150 4.4330 1.0780 ;
        RECT 1.9510 1.0780 4.4330 1.1280 ;
        RECT 1.9510 0.6700 2.0010 1.0780 ;
        RECT 2.2550 0.6700 2.3050 1.0780 ;
        RECT 3.1670 0.6700 3.2170 1.0780 ;
        RECT 3.4710 0.6700 3.5210 1.0780 ;
        RECT 3.7750 0.6700 3.8250 1.0780 ;
        RECT 4.0790 0.6700 4.1290 1.0780 ;
        RECT 2.5590 0.6700 2.6090 1.0780 ;
        RECT 2.8630 0.6700 2.9130 1.0780 ;
        RECT 4.3830 1.1280 4.4330 1.3140 ;
        RECT 0.8850 1.3140 4.4330 1.3640 ;
        RECT 1.1910 0.8540 1.2410 1.3140 ;
        RECT 1.4950 0.8540 1.5450 1.3140 ;
        RECT 0.8870 0.6710 0.9370 1.3140 ;
    END
  END VDDG

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4030 1.4440 1.6370 1.4940 ;
        RECT 1.4650 1.4940 1.5750 1.5750 ;
    END
    ANTENNAGATEAREA 0.0264 ;
  END D

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 5.3260 1.7020 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 5.3200 0.0300 ;
        RECT 1.1910 0.0300 1.2410 0.3000 ;
        RECT 1.9510 0.0300 2.0010 0.3510 ;
        RECT 2.5590 0.0300 2.6090 0.3510 ;
        RECT 2.8630 0.0300 2.9130 0.3510 ;
        RECT 3.4710 0.0300 3.5210 0.3510 ;
        RECT 3.1670 0.0300 3.2170 0.3510 ;
        RECT 4.0790 0.0300 4.1290 0.3510 ;
        RECT 3.7750 0.0300 3.8250 0.3510 ;
        RECT 2.2550 0.0300 2.3050 0.3510 ;
        RECT 0.8870 0.0300 0.9370 0.3260 ;
    END
  END VSS

  PIN ISO
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7950 0.4060 0.9670 0.4560 ;
        RECT 0.8570 0.4560 0.9670 0.4860 ;
        RECT 0.8570 0.3760 0.9670 0.4060 ;
    END
    ANTENNAGATEAREA 0.0186 ;
  END ISO
  OBS
    LAYER NWELL ;
      RECT 0.6540 0.4530 4.6870 1.0830 ;
      RECT -0.0910 1.5430 5.4410 1.7730 ;
      RECT -0.0910 0.6790 0.1940 1.5430 ;
      RECT 5.1470 0.6790 5.4410 1.5430 ;
    LAYER M1 ;
      RECT 0.7350 1.4290 1.3330 1.4790 ;
      RECT 0.7350 0.5710 0.7850 1.4290 ;
      RECT 0.6950 0.5210 0.7850 0.5710 ;
      RECT 0.6950 0.2890 0.7850 0.3390 ;
      RECT 0.7350 0.1210 0.7850 0.2890 ;
      RECT 0.6950 0.3390 0.7450 0.5210 ;
      RECT 1.3430 0.0880 1.6970 0.1380 ;
      RECT 1.6470 0.1380 1.6970 0.3000 ;
      RECT 1.3430 0.1380 1.3930 0.3500 ;
      RECT 1.0390 0.3500 1.3930 0.4000 ;
      RECT 1.0390 0.1260 1.0890 0.3500 ;
      RECT 1.6470 1.2140 4.2210 1.2640 ;
      RECT 1.0390 0.7670 1.0890 1.0180 ;
      RECT 1.3430 0.7670 1.3930 1.0280 ;
      RECT 1.6470 0.7670 1.6970 1.2140 ;
      RECT 1.0390 0.7170 1.6970 0.7670 ;
      RECT 1.4950 0.1980 1.5450 0.7170 ;
    LAYER PO ;
      RECT 3.1010 0.0710 3.1310 1.6040 ;
      RECT 3.2530 0.0710 3.2830 1.6030 ;
      RECT 3.4050 0.0710 3.4350 1.6100 ;
      RECT 3.5570 0.0700 3.5870 1.6030 ;
      RECT 3.7090 0.0710 3.7390 1.6040 ;
      RECT 3.8610 0.0710 3.8910 1.6040 ;
      RECT 4.0130 0.0710 4.0430 1.6030 ;
      RECT 4.1650 0.0710 4.1950 1.6100 ;
      RECT 1.4290 0.0710 1.4590 1.6030 ;
      RECT 1.5810 0.0710 1.6110 1.6040 ;
      RECT 2.4930 0.0710 2.5230 1.6040 ;
      RECT 0.8210 0.0710 0.8510 1.6030 ;
      RECT 0.9730 0.0710 1.0030 1.6030 ;
      RECT 0.6690 0.0710 0.6990 1.6030 ;
      RECT 2.0370 0.0710 2.0670 1.6100 ;
      RECT 0.5170 0.0710 0.5470 1.6040 ;
      RECT 2.7970 0.0710 2.8270 1.6100 ;
      RECT 0.3650 0.0710 0.3950 1.6030 ;
      RECT 2.6450 0.0710 2.6750 1.6030 ;
      RECT 1.1250 0.0710 1.1550 1.6030 ;
      RECT 1.7330 0.0720 1.7630 1.6040 ;
      RECT 2.1890 0.0700 2.2190 1.6030 ;
      RECT 1.2770 0.0710 1.3070 1.6040 ;
      RECT 1.8850 0.0710 1.9150 1.6030 ;
      RECT 2.3410 0.0710 2.3710 1.6040 ;
      RECT 2.9490 0.0710 2.9790 1.6100 ;
      RECT 4.7730 0.0710 4.8030 1.6100 ;
      RECT 4.6210 0.0710 4.6510 1.6100 ;
      RECT 4.4690 0.0710 4.4990 1.6030 ;
      RECT 4.3170 0.0710 4.3470 1.6040 ;
  END
END ISOLANDAOX8_LVT

MACRO ISOLANDX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.52 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.5200 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.2990 ;
        RECT 0.5830 0.0300 0.6330 0.4790 ;
        RECT 1.0390 0.0300 1.0890 0.5030 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.5200 1.7020 ;
        RECT 0.2790 1.1860 0.3290 1.6420 ;
        RECT 0.7350 1.1950 0.7850 1.6420 ;
        RECT 1.0390 0.8180 1.0890 1.6420 ;
    END
  END VDD

  PIN ISO
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2460 0.5830 0.4210 0.6330 ;
        RECT 0.2460 0.5530 0.3590 0.5830 ;
        RECT 0.2460 0.6330 0.3590 0.6630 ;
    END
    ANTENNAGATEAREA 0.0186 ;
  END ISO

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 0.8570 0.8150 0.8870 ;
        RECT 0.7050 0.8870 0.8770 0.9370 ;
        RECT 0.7050 0.9370 0.8150 0.9670 ;
    END
    ANTENNAGATEAREA 0.0234 ;
  END D

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1910 0.1170 1.2410 0.5470 ;
        RECT 1.1910 0.5470 1.3490 0.5530 ;
        RECT 1.1910 0.5530 1.4230 0.5970 ;
        RECT 1.2780 0.5970 1.4230 0.6630 ;
        RECT 1.2780 0.6630 1.3280 0.7580 ;
        RECT 1.1910 0.7580 1.3280 0.8080 ;
        RECT 1.1910 0.8080 1.2410 1.5590 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q
  OBS
    LAYER NWELL ;
      RECT -0.0910 0.6790 1.6350 1.7730 ;
    LAYER M1 ;
      RECT 0.4710 0.6970 0.7250 0.7470 ;
      RECT 0.4710 0.7470 0.5210 0.8590 ;
      RECT 0.4310 0.4580 0.5210 0.5080 ;
      RECT 0.4310 0.8590 0.5210 0.9090 ;
      RECT 0.4310 0.1170 0.4810 0.4580 ;
      RECT 0.4310 0.9090 0.4810 1.5590 ;
      RECT 0.4710 0.5080 0.5210 0.6970 ;
      RECT 0.8870 0.6560 1.1810 0.7060 ;
      RECT 0.8870 0.1060 0.9370 0.6560 ;
      RECT 0.9380 0.7060 0.9880 1.0930 ;
      RECT 0.5830 1.0930 0.9880 1.1430 ;
      RECT 0.8870 1.1430 0.9370 1.5680 ;
      RECT 0.5830 1.1430 0.6330 1.5680 ;
    LAYER PO ;
      RECT 0.3650 0.0670 0.3950 1.6050 ;
      RECT 0.2130 0.0660 0.2430 1.6030 ;
      RECT 0.5170 0.0670 0.5470 1.6030 ;
      RECT 0.9730 0.0660 1.0030 1.6030 ;
      RECT 1.1250 0.0670 1.1550 1.6050 ;
      RECT 1.4290 0.0670 1.4590 1.6030 ;
      RECT 1.2770 0.0670 1.3070 1.6030 ;
      RECT 0.0610 0.0660 0.0910 1.6030 ;
      RECT 0.8210 0.0660 0.8510 1.6030 ;
      RECT 0.6690 0.0660 0.6990 1.6030 ;
  END
END ISOLANDX1_LVT

MACRO ISOLANDX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.672 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN ISO
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2460 0.5830 0.4210 0.6330 ;
        RECT 0.2460 0.5530 0.3590 0.5830 ;
        RECT 0.2460 0.6330 0.3590 0.6630 ;
    END
    ANTENNAGATEAREA 0.0186 ;
  END ISO

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.6720 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.3030 ;
        RECT 0.5830 0.0300 0.6330 0.4790 ;
        RECT 1.1910 0.0300 1.2410 0.3980 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.6720 1.7020 ;
        RECT 0.2790 1.1860 0.3290 1.6420 ;
        RECT 0.7350 1.1950 0.7850 1.6420 ;
        RECT 1.1910 0.8080 1.2410 1.6420 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 0.7050 0.8150 0.7350 ;
        RECT 0.7050 0.7350 0.8770 0.7850 ;
        RECT 0.7050 0.7850 0.8150 0.8150 ;
    END
    ANTENNAGATEAREA 0.0234 ;
  END D

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0390 0.5030 1.4850 0.5530 ;
        RECT 1.4350 0.5530 1.5750 0.6630 ;
        RECT 1.3430 0.1300 1.3930 0.5030 ;
        RECT 1.0390 0.1300 1.0890 0.5030 ;
        RECT 1.4350 0.6630 1.4850 0.7080 ;
        RECT 1.0390 0.7080 1.4850 0.7580 ;
        RECT 1.0390 0.7580 1.0890 1.5440 ;
        RECT 1.3430 0.7580 1.3930 1.5440 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END Q
  OBS
    LAYER NWELL ;
      RECT -0.0910 0.6790 1.7870 1.7730 ;
    LAYER M1 ;
      RECT 0.4710 0.5960 0.7250 0.6460 ;
      RECT 0.4310 0.8590 0.5220 0.9090 ;
      RECT 0.4310 0.4580 0.5220 0.5080 ;
      RECT 0.4310 0.9090 0.4810 1.5590 ;
      RECT 0.4310 0.1170 0.4810 0.4580 ;
      RECT 0.4710 0.6460 0.5210 0.8590 ;
      RECT 0.4710 0.5080 0.5210 0.5960 ;
      RECT 0.9270 0.6080 1.3330 0.6580 ;
      RECT 0.9270 0.5740 0.9770 0.6080 ;
      RECT 0.6080 0.9390 0.9770 0.9400 ;
      RECT 0.8870 0.5240 0.9770 0.5740 ;
      RECT 0.5830 0.9400 0.9770 0.9890 ;
      RECT 0.8870 0.1210 0.9370 0.5240 ;
      RECT 0.8870 0.9890 0.9370 1.5530 ;
      RECT 0.9270 0.6580 0.9770 0.9390 ;
      RECT 0.5830 0.9890 0.6330 1.5530 ;
    LAYER PO ;
      RECT 0.0610 0.0710 0.0910 1.6030 ;
      RECT 0.2130 0.0710 0.2430 1.6030 ;
      RECT 0.3650 0.0710 0.3950 1.6040 ;
      RECT 1.5810 0.0720 1.6110 1.6100 ;
      RECT 0.5170 0.0710 0.5470 1.6030 ;
      RECT 0.8210 0.0710 0.8510 1.6030 ;
      RECT 0.6690 0.0710 0.6990 1.6030 ;
      RECT 0.9730 0.0710 1.0030 1.6030 ;
      RECT 1.1250 0.0720 1.1550 1.6040 ;
      RECT 1.4290 0.0720 1.4590 1.6030 ;
      RECT 1.2770 0.0720 1.3070 1.6040 ;
  END
END ISOLANDX2_LVT

MACRO ISOLANDX4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.976 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN ISO
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2460 0.5830 0.4210 0.6330 ;
        RECT 0.2460 0.5530 0.3590 0.5830 ;
        RECT 0.2460 0.6330 0.3590 0.6630 ;
    END
    ANTENNAGATEAREA 0.0186 ;
  END ISO

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7320 0.5530 1.8790 0.6630 ;
        RECT 1.7320 0.5330 1.7820 0.5530 ;
        RECT 1.7320 0.6630 1.7820 0.6930 ;
        RECT 1.0390 0.4830 1.7820 0.5330 ;
        RECT 1.0390 0.6930 1.7820 0.7430 ;
        RECT 1.0390 0.1150 1.0890 0.4830 ;
        RECT 1.3430 0.1150 1.3930 0.4830 ;
        RECT 1.6470 0.1150 1.6970 0.4830 ;
        RECT 1.0390 0.7430 1.0890 1.5440 ;
        RECT 1.3430 0.7430 1.3930 1.5440 ;
        RECT 1.6470 0.7430 1.6970 1.5440 ;
    END
    ANTENNADIFFAREA 0.3972 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.9760 1.7020 ;
        RECT 0.2790 1.1860 0.3290 1.6420 ;
        RECT 1.1910 0.8180 1.2410 1.6420 ;
        RECT 1.4950 0.8180 1.5450 1.6420 ;
        RECT 0.7350 1.2880 0.7850 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.9760 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.3030 ;
        RECT 1.1910 0.0300 1.2410 0.4130 ;
        RECT 0.5830 0.0300 0.6330 0.4800 ;
        RECT 1.4950 0.0300 1.5450 0.4130 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 0.7050 0.8150 0.7350 ;
        RECT 0.7050 0.7350 0.8770 0.7850 ;
        RECT 0.7050 0.7850 0.8150 0.8150 ;
    END
    ANTENNAGATEAREA 0.0228 ;
  END D
  OBS
    LAYER NWELL ;
      RECT -0.0910 0.6790 2.0910 1.7730 ;
    LAYER M1 ;
      RECT 0.4710 0.5960 0.7250 0.6460 ;
      RECT 0.4310 0.8590 0.5220 0.9090 ;
      RECT 0.4310 0.4580 0.5220 0.5080 ;
      RECT 0.4310 0.9090 0.4810 1.5590 ;
      RECT 0.4310 0.1170 0.4810 0.4580 ;
      RECT 0.4710 0.6460 0.5210 0.8590 ;
      RECT 0.4710 0.5080 0.5210 0.5960 ;
      RECT 0.8870 0.5910 1.6370 0.6410 ;
      RECT 0.8870 0.1220 0.9370 0.5910 ;
      RECT 0.9280 0.6410 0.9780 0.8670 ;
      RECT 0.5830 0.8670 0.9780 0.9170 ;
      RECT 0.8870 0.9170 0.9370 1.5540 ;
      RECT 0.5830 0.9170 0.6330 1.5540 ;
    LAYER PO ;
      RECT 0.0610 0.0710 0.0910 1.6030 ;
      RECT 0.2130 0.0710 0.2430 1.6030 ;
      RECT 0.3650 0.0710 0.3950 1.6040 ;
      RECT 1.2770 0.0720 1.3070 1.6040 ;
      RECT 1.4290 0.0720 1.4590 1.6040 ;
      RECT 1.5810 0.0720 1.6110 1.6040 ;
      RECT 1.8850 0.0720 1.9150 1.6040 ;
      RECT 1.7330 0.0720 1.7630 1.6040 ;
      RECT 1.1250 0.0720 1.1550 1.6040 ;
      RECT 0.9730 0.0710 1.0030 1.6040 ;
      RECT 0.6690 0.0710 0.6990 1.6040 ;
      RECT 0.8210 0.0710 0.8510 1.6040 ;
      RECT 0.5170 0.0710 0.5470 1.6040 ;
  END
END ISOLANDX4_LVT

MACRO ISOLANDX8_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.584 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 0.7050 0.8150 0.7350 ;
        RECT 0.7050 0.7350 0.8770 0.7850 ;
        RECT 0.7050 0.7850 0.8150 0.8150 ;
    END
    ANTENNAGATEAREA 0.0234 ;
  END D

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.5840 0.0300 ;
        RECT 1.7990 0.0300 1.8490 0.4130 ;
        RECT 2.1030 0.0300 2.1530 0.4130 ;
        RECT 0.2790 0.0300 0.3290 0.3030 ;
        RECT 1.4950 0.0300 1.5450 0.4130 ;
        RECT 1.1910 0.0300 1.2410 0.4130 ;
        RECT 0.5830 0.0300 0.6330 0.4800 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.5840 1.7020 ;
        RECT 1.7990 0.8180 1.8490 1.6420 ;
        RECT 2.1030 0.8180 2.1530 1.6420 ;
        RECT 0.2790 1.1860 0.3290 1.6420 ;
        RECT 0.7350 1.1960 0.7850 1.6420 ;
        RECT 1.4950 0.8180 1.5450 1.6420 ;
        RECT 1.1910 0.8180 1.2410 1.6420 ;
    END
  END VDD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3750 0.5330 2.4250 0.5530 ;
        RECT 2.3750 0.5530 2.4870 0.6630 ;
        RECT 1.0390 0.4830 2.4250 0.5330 ;
        RECT 2.3750 0.6630 2.4250 0.7030 ;
        RECT 1.9510 0.1150 2.0010 0.4830 ;
        RECT 2.2550 0.1150 2.3050 0.4830 ;
        RECT 1.6470 0.1150 1.6970 0.4830 ;
        RECT 1.3430 0.1150 1.3930 0.4830 ;
        RECT 1.0390 0.1150 1.0890 0.4830 ;
        RECT 1.0390 0.7030 2.4250 0.7530 ;
        RECT 1.9510 0.7530 2.0010 1.5440 ;
        RECT 2.2550 0.7530 2.3050 1.5440 ;
        RECT 1.6470 0.7530 1.6970 1.5440 ;
        RECT 1.3430 0.7530 1.3930 1.5440 ;
        RECT 1.0390 0.7530 1.0890 1.5440 ;
    END
    ANTENNADIFFAREA 0.6952 ;
  END Q

  PIN ISO
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2460 0.5530 0.3590 0.5830 ;
        RECT 0.2460 0.5830 0.4210 0.6330 ;
        RECT 0.2460 0.6330 0.3590 0.6630 ;
    END
    ANTENNAGATEAREA 0.0186 ;
  END ISO
  OBS
    LAYER NWELL ;
      RECT -0.0910 0.6790 2.6750 1.7730 ;
    LAYER M1 ;
      RECT 0.4310 0.8590 0.5220 0.9090 ;
      RECT 0.4310 0.4580 0.5220 0.5080 ;
      RECT 0.4310 0.9090 0.4810 1.5590 ;
      RECT 0.4310 0.1170 0.4810 0.4580 ;
      RECT 0.4710 0.5960 0.7250 0.6460 ;
      RECT 0.4710 0.6460 0.5210 0.8590 ;
      RECT 0.4710 0.5080 0.5210 0.5960 ;
      RECT 0.8870 0.5910 2.3250 0.6410 ;
      RECT 0.5830 0.9170 0.6330 1.5540 ;
      RECT 0.8870 0.1220 0.9370 0.5910 ;
      RECT 0.5830 0.8670 0.9770 0.9170 ;
      RECT 0.8870 0.9170 0.9370 1.5540 ;
      RECT 0.9270 0.6410 0.9770 0.8670 ;
    LAYER PO ;
      RECT 2.4930 0.0720 2.5230 1.6040 ;
      RECT 2.3410 0.0720 2.3710 1.6040 ;
      RECT 2.1890 0.0720 2.2190 1.6040 ;
      RECT 2.0370 0.0720 2.0670 1.6040 ;
      RECT 0.5170 0.0710 0.5470 1.6040 ;
      RECT 0.8210 0.0710 0.8510 1.6040 ;
      RECT 0.6690 0.0710 0.6990 1.6040 ;
      RECT 0.9730 0.0710 1.0030 1.6040 ;
      RECT 1.1250 0.0720 1.1550 1.6040 ;
      RECT 1.7330 0.0720 1.7630 1.6040 ;
      RECT 1.8850 0.0720 1.9150 1.6040 ;
      RECT 1.5810 0.0720 1.6110 1.6040 ;
      RECT 1.4290 0.0720 1.4590 1.6040 ;
      RECT 1.2770 0.0720 1.3070 1.6040 ;
      RECT 0.3650 0.0710 0.3950 1.6040 ;
      RECT 0.2130 0.0710 0.2430 1.6030 ;
      RECT 0.0610 0.0710 0.0910 1.6030 ;
  END
END ISOLANDX8_LVT

MACRO ISOLORAOX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.496 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 2.5290 0.7050 2.6390 0.8150 ;
        RECT 2.5590 0.6830 2.6090 0.7050 ;
        RECT 2.5590 0.8150 2.6090 1.0780 ;
        RECT 1.7990 1.0780 2.6090 1.1280 ;
        RECT 1.7990 0.8540 1.8490 1.0780 ;
        RECT 2.2550 0.7620 2.3050 1.0780 ;
    END
  END VDDG

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.7350 0.5110 0.7850 ;
        RECT 0.4010 0.7050 0.5110 0.7350 ;
        RECT 0.4010 0.7850 0.5110 0.8150 ;
    END
    ANTENNAGATEAREA 0.0186 ;
  END D

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.4960 1.7020 ;
        RECT 0.4310 1.1960 0.4810 1.6420 ;
    END
  END VDD

  PIN ISO
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7070 1.3430 1.9410 1.3930 ;
        RECT 1.7690 1.3930 1.8790 1.4230 ;
        RECT 1.7690 1.3130 1.8790 1.3430 ;
    END
    ANTENNAGATEAREA 0.0312 ;
  END ISO

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.4960 0.0300 ;
        RECT 1.6470 0.0300 1.6970 0.2130 ;
        RECT 1.3430 0.0300 1.3930 0.2130 ;
        RECT 1.9510 0.0300 2.0010 0.2130 ;
        RECT 2.2550 0.0300 2.3050 0.2130 ;
        RECT 0.4310 0.0300 0.4810 0.2950 ;
    END
  END VSS

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5290 0.4010 2.6400 0.4910 ;
        RECT 2.4070 0.4910 2.6400 0.5410 ;
        RECT 2.5490 0.3130 2.5990 0.4010 ;
        RECT 2.4070 0.5410 2.4570 0.6620 ;
        RECT 2.1030 0.2630 2.5990 0.3130 ;
        RECT 2.1030 0.6620 2.4570 0.7120 ;
        RECT 2.4070 0.1310 2.4570 0.2630 ;
        RECT 2.1030 0.1310 2.1530 0.2630 ;
        RECT 2.1030 0.7120 2.1530 1.0280 ;
        RECT 2.4070 0.7120 2.4570 1.0280 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q
  OBS
    LAYER NWELL ;
      RECT -0.0910 1.5430 3.6110 1.7730 ;
      RECT -0.0910 0.6790 0.7190 1.5430 ;
      RECT 3.3230 0.6790 3.6110 1.5430 ;
      RECT 1.1790 0.4530 2.8630 1.0830 ;
    LAYER M1 ;
      RECT 0.7950 1.3430 1.6370 1.3930 ;
      RECT 0.7950 0.7480 0.8450 1.3430 ;
      RECT 0.6230 0.6980 0.8450 0.7480 ;
      RECT 0.7950 0.6970 0.8450 0.6980 ;
      RECT 0.6230 0.5730 0.6730 0.6980 ;
      RECT 0.6230 0.7480 0.6730 1.1200 ;
      RECT 0.5830 0.5230 0.6730 0.5730 ;
      RECT 0.5830 1.1200 0.6730 1.1700 ;
      RECT 0.5830 0.1140 0.6330 0.5230 ;
      RECT 0.5830 1.1700 0.6330 1.5610 ;
      RECT 0.2390 0.9810 0.5730 1.0310 ;
      RECT 0.2390 1.0310 0.2890 1.0960 ;
      RECT 0.2390 1.0960 0.3290 1.1700 ;
      RECT 0.2390 0.5040 0.3290 0.5540 ;
      RECT 0.2790 1.1700 0.3290 1.5540 ;
      RECT 0.2790 0.1210 0.3290 0.5040 ;
      RECT 0.2390 0.5540 0.2890 0.9810 ;
      RECT 1.6470 0.6700 2.0010 0.7200 ;
      RECT 1.9510 0.7200 2.0010 1.0280 ;
      RECT 1.6470 0.7200 1.6970 1.0780 ;
      RECT 1.3430 1.0780 1.6970 1.1280 ;
      RECT 1.3430 0.7620 1.3930 1.0780 ;
      RECT 1.4950 0.3770 2.3970 0.4270 ;
      RECT 1.4950 0.4270 1.5450 1.0280 ;
      RECT 1.4950 0.1260 1.5450 0.3770 ;
      RECT 1.7990 0.1310 1.8490 0.3770 ;
    LAYER PO ;
      RECT 0.0610 0.0710 0.0910 1.6040 ;
      RECT 0.5170 0.0710 0.5470 1.6040 ;
      RECT 0.3650 0.0710 0.3950 1.6040 ;
      RECT 0.6690 0.0710 0.6990 1.6040 ;
      RECT 0.8210 0.0710 0.8510 1.6040 ;
      RECT 2.0370 0.0720 2.0670 1.6040 ;
      RECT 0.9730 0.0710 1.0030 1.6040 ;
      RECT 1.2770 0.0710 1.3070 1.6040 ;
      RECT 1.1250 0.0710 1.1550 1.6040 ;
      RECT 2.4930 0.0710 2.5230 1.6040 ;
      RECT 1.4290 0.0710 1.4590 1.6040 ;
      RECT 1.5810 0.0710 1.6110 1.6040 ;
      RECT 1.8850 0.0710 1.9150 1.6040 ;
      RECT 1.7330 0.0710 1.7630 1.6040 ;
      RECT 2.1890 0.0710 2.2190 1.6040 ;
      RECT 2.3410 0.0710 2.3710 1.6040 ;
      RECT 2.6450 0.0720 2.6750 1.6040 ;
      RECT 2.7970 0.0720 2.8270 1.6040 ;
      RECT 0.2130 0.0710 0.2430 1.6040 ;
  END
END ISOLORAOX1_LVT

MACRO ISOLORAOX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.8330 0.4010 2.9440 0.4780 ;
        RECT 2.8530 0.3130 2.9030 0.4010 ;
        RECT 2.7110 0.4780 2.9440 0.5080 ;
        RECT 2.1030 0.2630 2.9030 0.3130 ;
        RECT 2.1240 0.5080 2.9440 0.5090 ;
        RECT 2.7110 0.1310 2.7610 0.2630 ;
        RECT 2.1030 0.1310 2.1530 0.2630 ;
        RECT 2.4070 0.1310 2.4570 0.2630 ;
        RECT 2.1030 0.5090 2.9440 0.5280 ;
        RECT 2.1030 0.5280 2.7610 0.5580 ;
        RECT 2.1030 0.5580 2.1530 1.0280 ;
        RECT 2.4070 0.5580 2.4570 1.0280 ;
        RECT 2.7110 0.5580 2.7610 1.0280 ;
    END
    ANTENNADIFFAREA 0.1988 ;
  END Q

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.8000 0.0300 ;
        RECT 2.5590 0.0300 2.6090 0.2130 ;
        RECT 2.2550 0.0300 2.3050 0.2130 ;
        RECT 0.4310 0.0300 0.4810 0.2950 ;
        RECT 1.6470 0.0300 1.6970 0.2130 ;
        RECT 1.9510 0.0300 2.0010 0.2130 ;
        RECT 1.3430 0.0300 1.3930 0.2130 ;
    END
  END VSS

  PIN ISO
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7070 1.3430 1.9410 1.3930 ;
        RECT 1.7690 1.3930 1.8790 1.4230 ;
        RECT 1.7690 1.3130 1.8790 1.3430 ;
    END
    ANTENNAGATEAREA 0.0312 ;
  END ISO

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.8000 1.7020 ;
        RECT 0.4310 1.1960 0.4810 1.6420 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.7350 0.5110 0.7850 ;
        RECT 0.4010 0.7850 0.5110 0.8150 ;
        RECT 0.4010 0.7050 0.5110 0.7350 ;
    END
    ANTENNAGATEAREA 0.0186 ;
  END D

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 2.8330 0.7050 2.9430 0.8150 ;
        RECT 2.8630 0.6830 2.9130 0.7050 ;
        RECT 2.8630 0.8150 2.9130 1.0780 ;
        RECT 1.7990 1.0780 2.9130 1.1280 ;
        RECT 1.7990 0.6700 1.8490 1.0780 ;
        RECT 2.5590 0.6700 2.6090 1.0780 ;
        RECT 2.2550 0.6700 2.3050 1.0780 ;
    END
  END VDDG
  OBS
    LAYER NWELL ;
      RECT -0.0910 1.5430 3.9150 1.7730 ;
      RECT -0.0910 0.6790 0.7190 1.5430 ;
      RECT 3.6270 0.6790 3.9150 1.5430 ;
      RECT 1.1790 0.4530 3.1670 1.0830 ;
    LAYER M1 ;
      RECT 0.2390 0.9810 0.5730 1.0310 ;
      RECT 0.2390 1.0310 0.2890 1.0960 ;
      RECT 0.2390 0.5040 0.3290 0.5540 ;
      RECT 0.2390 1.0960 0.3290 1.1700 ;
      RECT 0.2790 0.1210 0.3290 0.5040 ;
      RECT 0.2790 1.1700 0.3290 1.5540 ;
      RECT 0.2390 0.5540 0.2890 0.9810 ;
      RECT 0.7950 1.3430 1.6370 1.3930 ;
      RECT 0.7950 0.7480 0.8450 1.3430 ;
      RECT 0.6230 0.6980 0.8450 0.7480 ;
      RECT 0.7950 0.6970 0.8450 0.6980 ;
      RECT 0.6230 0.7480 0.6730 1.1200 ;
      RECT 0.6230 0.5740 0.6730 0.6980 ;
      RECT 0.5830 1.1200 0.6730 1.1700 ;
      RECT 0.5830 0.5240 0.6730 0.5740 ;
      RECT 0.5830 1.1700 0.6330 1.5610 ;
      RECT 0.5830 0.1140 0.6330 0.5240 ;
      RECT 1.6470 0.5440 2.0010 0.5940 ;
      RECT 1.9510 0.5940 2.0010 1.0280 ;
      RECT 1.6470 0.5940 1.6970 1.0780 ;
      RECT 1.3430 1.0780 1.6970 1.1280 ;
      RECT 1.3430 0.6700 1.3930 1.0780 ;
      RECT 1.4950 0.3770 2.7010 0.4270 ;
      RECT 1.4950 0.4270 1.5450 1.0280 ;
      RECT 1.4950 0.1260 1.5450 0.3770 ;
      RECT 1.7990 0.1310 1.8490 0.3770 ;
    LAYER PO ;
      RECT 2.4930 0.0710 2.5230 1.6040 ;
      RECT 1.4290 0.0710 1.4590 1.6040 ;
      RECT 1.5810 0.0710 1.6110 1.6040 ;
      RECT 1.8850 0.0710 1.9150 1.6040 ;
      RECT 1.7330 0.0710 1.7630 1.6040 ;
      RECT 2.1890 0.0710 2.2190 1.6040 ;
      RECT 3.2530 0.0710 3.2830 1.6040 ;
      RECT 3.5570 0.0710 3.5870 1.6040 ;
      RECT 0.2130 0.0710 0.2430 1.6040 ;
      RECT 2.9490 0.0710 2.9790 1.6040 ;
      RECT 2.7970 0.0710 2.8270 1.6040 ;
      RECT 2.6450 0.0710 2.6750 1.6040 ;
      RECT 2.3410 0.0710 2.3710 1.6040 ;
      RECT 3.1010 0.0710 3.1310 1.6040 ;
      RECT 0.3650 0.0710 0.3950 1.6040 ;
      RECT 0.5170 0.0710 0.5470 1.6040 ;
      RECT 0.0610 0.0710 0.0910 1.6040 ;
      RECT 3.4050 0.0710 3.4350 1.6040 ;
      RECT 1.1250 0.0710 1.1550 1.6040 ;
      RECT 1.2770 0.0710 1.3070 1.6040 ;
      RECT 0.9730 0.0710 1.0030 1.6040 ;
      RECT 2.0370 0.0720 2.0670 1.6040 ;
      RECT 0.8210 0.0710 0.8510 1.6040 ;
      RECT 0.6690 0.0710 0.6990 1.6040 ;
  END
END ISOLORAOX2_LVT

MACRO HEADX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.128 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDDG
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.6660 1.0090 0.8560 1.1190 ;
        RECT 0.7300 1.1190 0.7900 1.1650 ;
        RECT 0.7300 0.8810 0.7900 1.0090 ;
        RECT 0.7300 0.8560 1.2410 0.8810 ;
        RECT 0.7350 0.8310 1.2410 0.8560 ;
        RECT 1.1910 0.8810 1.2410 1.5610 ;
    END
  END VDDG

  PIN VDD
    DIRECTION OUTPUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.1280 1.7020 ;
        RECT 1.0390 1.0150 1.0890 1.6420 ;
        RECT 1.3430 1.0150 1.3930 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.1280 0.0300 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 2.1280 3.3740 ;
    END
  END VSS

  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0990 0.6700 1.3330 0.7300 ;
        RECT 1.1200 0.5530 1.3100 0.6700 ;
    END
  END SLEEP
  OBS
    LAYER NWELL ;
      RECT 0.5710 0.6790 1.5490 2.6650 ;
    LAYER PO ;
      RECT 0.0610 0.1230 0.0910 1.6210 ;
      RECT 0.2130 0.1230 0.2430 1.6210 ;
      RECT 0.3650 0.1230 0.3950 1.6210 ;
      RECT 0.5170 0.1230 0.5470 1.6210 ;
      RECT 1.5810 0.1230 1.6110 1.6210 ;
      RECT 2.0370 0.1230 2.0670 1.6210 ;
      RECT 1.8850 0.1230 1.9150 1.6210 ;
      RECT 1.7330 0.1230 1.7630 1.6210 ;
      RECT 0.0610 1.7670 0.0910 3.2650 ;
      RECT 0.2130 1.7670 0.2430 3.2650 ;
      RECT 0.3650 1.7670 0.3950 3.2650 ;
      RECT 0.5170 1.7670 0.5470 3.2650 ;
      RECT 1.5810 1.7670 1.6110 3.2650 ;
      RECT 2.0370 1.7670 2.0670 3.2650 ;
      RECT 1.8850 1.7670 1.9150 3.2650 ;
      RECT 1.7330 1.7670 1.7630 3.2650 ;
      RECT 1.1250 1.7670 1.1550 3.2650 ;
      RECT 1.2770 1.7670 1.3070 3.2650 ;
      RECT 1.4290 1.7670 1.4590 3.2650 ;
      RECT 0.9730 1.7670 1.0030 3.2650 ;
      RECT 0.8210 1.7670 0.8510 3.2650 ;
      RECT 0.6690 1.7670 0.6990 3.2650 ;
      RECT 0.6690 0.1230 0.6990 1.6210 ;
      RECT 0.8210 0.1230 0.8510 1.6210 ;
      RECT 0.9730 0.1230 1.0030 1.6210 ;
      RECT 1.4290 0.1230 1.4590 1.6210 ;
      RECT 1.2770 0.1230 1.3070 1.6210 ;
      RECT 1.1250 0.1230 1.1550 1.6210 ;
  END
END HEADX2_LVT

MACRO HEADX32_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.688 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDDG
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.6660 1.0090 0.8560 1.1190 ;
        RECT 0.7300 1.1190 0.7900 1.1650 ;
        RECT 0.7300 0.8810 0.7900 1.0090 ;
        RECT 0.7300 0.8560 5.8010 0.8810 ;
        RECT 0.7350 0.8310 5.8010 0.8560 ;
        RECT 1.7990 0.8810 1.8490 1.5610 ;
        RECT 1.4950 0.8810 1.5450 1.5610 ;
        RECT 1.1910 0.8810 1.2410 1.5610 ;
        RECT 3.3190 0.8810 3.3690 1.5610 ;
        RECT 3.6230 0.8810 3.6730 1.5610 ;
        RECT 3.9270 0.8810 3.9770 1.5610 ;
        RECT 4.2310 0.8810 4.2810 1.5610 ;
        RECT 4.5350 0.8810 4.5850 1.5610 ;
        RECT 4.8390 0.8810 4.8890 1.5610 ;
        RECT 5.1430 0.8810 5.1930 1.5610 ;
        RECT 5.4470 0.8810 5.4970 1.5610 ;
        RECT 2.1030 0.8810 2.1530 1.5610 ;
        RECT 2.4070 0.8810 2.4570 1.5610 ;
        RECT 2.7110 0.8810 2.7610 1.5610 ;
        RECT 3.0150 0.8810 3.0650 1.5610 ;
        RECT 5.7510 0.8810 5.8010 1.5610 ;
    END
  END VDDG

  PIN VDD
    DIRECTION OUTPUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 6.6880 1.7020 ;
        RECT 5.9030 0.8330 5.9530 1.6420 ;
        RECT 5.5990 1.0170 5.6490 1.6420 ;
        RECT 5.2950 1.0170 5.3450 1.6420 ;
        RECT 4.9910 1.0170 5.0410 1.6420 ;
        RECT 4.6870 1.0170 4.7370 1.6420 ;
        RECT 4.3830 1.0170 4.4330 1.6420 ;
        RECT 4.0790 1.0170 4.1290 1.6420 ;
        RECT 3.7750 1.0170 3.8250 1.6420 ;
        RECT 3.4710 1.0170 3.5210 1.6420 ;
        RECT 3.1670 1.0170 3.2170 1.6420 ;
        RECT 2.8630 1.0170 2.9130 1.6420 ;
        RECT 2.5590 1.0170 2.6090 1.6420 ;
        RECT 2.2550 1.0170 2.3050 1.6420 ;
        RECT 1.9510 1.0170 2.0010 1.6420 ;
        RECT 1.0390 1.0170 1.0890 1.6420 ;
        RECT 1.6470 1.0170 1.6970 1.6420 ;
        RECT 1.3430 1.0170 1.3930 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 6.6880 0.0300 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 6.6880 3.3740 ;
    END
  END VSS

  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0990 0.6700 5.8930 0.7300 ;
        RECT 1.1200 0.5530 1.3100 0.6700 ;
    END
  END SLEEP
  OBS
    LAYER NWELL ;
      RECT 0.5710 0.6790 6.1090 2.6650 ;
    LAYER PO ;
      RECT 1.1250 1.7460 1.1550 3.2640 ;
      RECT 1.2770 1.7460 1.3070 3.2640 ;
      RECT 3.7090 1.7460 3.7390 3.2640 ;
      RECT 3.8610 1.7460 3.8910 3.2640 ;
      RECT 4.0130 1.7460 4.0430 3.2640 ;
      RECT 4.1650 1.7460 4.1950 3.2640 ;
      RECT 4.3170 1.7460 4.3470 3.2640 ;
      RECT 4.4690 1.7460 4.4990 3.2640 ;
      RECT 4.6210 1.7460 4.6510 3.2640 ;
      RECT 4.7730 1.7460 4.8030 3.2640 ;
      RECT 4.9250 1.7460 4.9550 3.2640 ;
      RECT 5.0770 1.7460 5.1070 3.2640 ;
      RECT 5.2290 1.7460 5.2590 3.2640 ;
      RECT 5.3810 1.7460 5.4110 3.2640 ;
      RECT 5.5330 1.7460 5.5630 3.2640 ;
      RECT 5.6850 1.7460 5.7150 3.2640 ;
      RECT 5.9890 1.7460 6.0190 3.2640 ;
      RECT 2.0370 1.7460 2.0670 3.2640 ;
      RECT 1.8850 1.7460 1.9150 3.2640 ;
      RECT 0.6690 1.7460 0.6990 3.2640 ;
      RECT 0.0610 0.1030 0.0910 1.6210 ;
      RECT 0.2130 0.1030 0.2430 1.6210 ;
      RECT 0.3650 0.1030 0.3950 1.6210 ;
      RECT 0.5170 0.1030 0.5470 1.6210 ;
      RECT 6.1410 0.1030 6.1710 1.6210 ;
      RECT 6.2930 0.1030 6.3230 1.6210 ;
      RECT 6.4450 0.1030 6.4750 1.6210 ;
      RECT 6.5970 0.1030 6.6270 1.6210 ;
      RECT 6.5970 1.7460 6.6270 3.2640 ;
      RECT 6.4450 1.7460 6.4750 3.2640 ;
      RECT 6.2930 1.7460 6.3230 3.2640 ;
      RECT 6.1410 1.7460 6.1710 3.2640 ;
      RECT 0.5170 1.7460 0.5470 3.2640 ;
      RECT 0.3650 1.7460 0.3950 3.2640 ;
      RECT 0.2130 1.7460 0.2430 3.2640 ;
      RECT 0.0610 1.7460 0.0910 3.2640 ;
      RECT 2.6450 1.7460 2.6750 3.2640 ;
      RECT 2.4930 1.7460 2.5230 3.2640 ;
      RECT 3.5570 1.7460 3.5870 3.2640 ;
      RECT 2.3410 1.7460 2.3710 3.2640 ;
      RECT 2.1890 1.7460 2.2190 3.2640 ;
      RECT 2.7970 1.7460 2.8270 3.2640 ;
      RECT 2.9490 1.7460 2.9790 3.2640 ;
      RECT 3.1010 1.7460 3.1310 3.2640 ;
      RECT 3.2530 1.7460 3.2830 3.2640 ;
      RECT 3.4050 1.7460 3.4350 3.2640 ;
      RECT 2.6450 0.1030 2.6750 1.6210 ;
      RECT 2.4930 0.1030 2.5230 1.6210 ;
      RECT 3.5570 0.1030 3.5870 1.6210 ;
      RECT 2.3410 0.1030 2.3710 1.6210 ;
      RECT 2.1890 0.1030 2.2190 1.6210 ;
      RECT 2.0370 0.1030 2.0670 1.6210 ;
      RECT 1.8850 0.1030 1.9150 1.6210 ;
      RECT 0.6690 0.1030 0.6990 1.6210 ;
      RECT 1.5810 0.1030 1.6110 1.6210 ;
      RECT 0.8210 0.1030 0.8510 1.6210 ;
      RECT 0.9730 0.1030 1.0030 1.6210 ;
      RECT 1.4290 0.1030 1.4590 1.6210 ;
      RECT 1.7330 0.1030 1.7630 1.6210 ;
      RECT 1.1250 0.1030 1.1550 1.6210 ;
      RECT 1.2770 0.1030 1.3070 1.6210 ;
      RECT 3.7090 0.1030 3.7390 1.6210 ;
      RECT 3.8610 0.1030 3.8910 1.6210 ;
      RECT 4.0130 0.1030 4.0430 1.6210 ;
      RECT 4.1650 0.1030 4.1950 1.6210 ;
      RECT 4.3170 0.1030 4.3470 1.6210 ;
      RECT 4.4690 0.1030 4.4990 1.6210 ;
      RECT 4.6210 0.1030 4.6510 1.6210 ;
      RECT 4.7730 0.1030 4.8030 1.6210 ;
      RECT 4.9250 0.1030 4.9550 1.6210 ;
      RECT 5.0770 0.1030 5.1070 1.6210 ;
      RECT 5.2290 0.1030 5.2590 1.6210 ;
      RECT 5.3810 0.1030 5.4110 1.6210 ;
      RECT 5.5330 0.1030 5.5630 1.6210 ;
      RECT 5.6850 0.1030 5.7150 1.6210 ;
      RECT 5.8370 0.1030 5.8670 1.6210 ;
      RECT 5.9890 0.1030 6.0190 1.6210 ;
      RECT 3.4050 0.1030 3.4350 1.6210 ;
      RECT 3.2530 0.1030 3.2830 1.6210 ;
      RECT 3.1010 0.1030 3.1310 1.6210 ;
      RECT 2.9490 0.1030 2.9790 1.6210 ;
      RECT 2.7970 0.1030 2.8270 1.6210 ;
      RECT 5.8370 1.7460 5.8670 3.2640 ;
      RECT 1.5810 1.7460 1.6110 3.2640 ;
      RECT 0.8210 1.7460 0.8510 3.2640 ;
      RECT 0.9730 1.7460 1.0030 3.2640 ;
      RECT 1.4290 1.7460 1.4590 3.2640 ;
      RECT 1.7330 1.7460 1.7630 3.2640 ;
  END
END HEADX32_LVT

MACRO HEADX4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.432 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDDG
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.6660 1.0090 0.8560 1.1190 ;
        RECT 0.7300 1.1190 0.7900 1.1650 ;
        RECT 0.7300 0.8810 0.7900 1.0090 ;
        RECT 0.7300 0.8560 1.5450 0.8810 ;
        RECT 0.7350 0.8310 1.5450 0.8560 ;
        RECT 1.1910 0.8810 1.2410 1.5610 ;
        RECT 1.4950 0.8810 1.5450 1.5610 ;
    END
  END VDDG

  PIN VDD
    DIRECTION OUTPUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.4320 1.7020 ;
        RECT 1.0390 1.0170 1.0890 1.6420 ;
        RECT 1.6470 0.8330 1.6970 1.6420 ;
        RECT 1.3430 1.0170 1.3930 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.4320 0.0300 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 2.4320 3.3740 ;
    END
  END VSS

  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0990 0.6700 1.6370 0.7300 ;
        RECT 1.1200 0.5530 1.3100 0.6700 ;
    END
  END SLEEP
  OBS
    LAYER NWELL ;
      RECT 0.5710 0.6790 1.8530 2.6650 ;
    LAYER PO ;
      RECT 0.5170 0.1130 0.5470 1.6210 ;
      RECT 0.3650 0.1130 0.3950 1.6210 ;
      RECT 0.2130 0.1130 0.2430 1.6210 ;
      RECT 0.0610 0.1130 0.0910 1.6210 ;
      RECT 1.8850 0.1130 1.9150 1.6210 ;
      RECT 2.3410 0.1130 2.3710 1.6210 ;
      RECT 2.0370 0.1130 2.0670 1.6210 ;
      RECT 2.1890 0.1130 2.2190 1.6210 ;
      RECT 0.0610 1.7580 0.0910 3.2660 ;
      RECT 0.2130 1.7580 0.2430 3.2660 ;
      RECT 0.3650 1.7580 0.3950 3.2660 ;
      RECT 0.5170 1.7580 0.5470 3.2660 ;
      RECT 1.8850 1.7580 1.9150 3.2660 ;
      RECT 2.3410 1.7580 2.3710 3.2660 ;
      RECT 2.0370 1.7580 2.0670 3.2660 ;
      RECT 2.1890 1.7580 2.2190 3.2660 ;
      RECT 1.2770 1.7580 1.3070 3.2660 ;
      RECT 1.1250 1.7580 1.1550 3.2660 ;
      RECT 1.7330 1.7580 1.7630 3.2660 ;
      RECT 1.4290 1.7580 1.4590 3.2660 ;
      RECT 0.9730 1.7580 1.0030 3.2660 ;
      RECT 0.8210 1.7580 0.8510 3.2660 ;
      RECT 1.5810 1.7580 1.6110 3.2660 ;
      RECT 0.6690 1.7580 0.6990 3.2660 ;
      RECT 0.6690 0.1130 0.6990 1.6210 ;
      RECT 1.5810 0.1130 1.6110 1.6210 ;
      RECT 0.8210 0.1130 0.8510 1.6210 ;
      RECT 0.9730 0.1130 1.0030 1.6210 ;
      RECT 1.4290 0.1130 1.4590 1.6210 ;
      RECT 1.7330 0.1130 1.7630 1.6210 ;
      RECT 1.1250 0.1130 1.1550 1.6210 ;
      RECT 1.2770 0.1130 1.3070 1.6210 ;
  END
END HEADX4_LVT

MACRO HEADX8_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.04 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDDG
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.6660 1.0090 0.8560 1.1190 ;
        RECT 0.7300 1.1190 0.7900 1.1650 ;
        RECT 0.7300 0.8810 0.7900 1.0090 ;
        RECT 0.7300 0.8560 2.1530 0.8810 ;
        RECT 0.7350 0.8310 2.1530 0.8560 ;
        RECT 1.7990 0.8810 1.8490 1.5610 ;
        RECT 1.4950 0.8810 1.5450 1.5610 ;
        RECT 1.1910 0.8810 1.2410 1.5610 ;
        RECT 2.1030 0.8810 2.1530 1.5610 ;
    END
  END VDDG

  PIN VDD
    DIRECTION OUTPUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.0400 1.7020 ;
        RECT 2.2550 0.8330 2.3050 1.6420 ;
        RECT 1.9510 1.0170 2.0010 1.6420 ;
        RECT 1.0390 1.0170 1.0890 1.6420 ;
        RECT 1.6470 1.0170 1.6970 1.6420 ;
        RECT 1.3430 1.0170 1.3930 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.0400 0.0300 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 3.0400 3.3740 ;
    END
  END VSS

  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0990 0.6700 2.2450 0.7300 ;
        RECT 1.1200 0.5530 1.3100 0.6700 ;
    END
  END SLEEP
  OBS
    LAYER NWELL ;
      RECT 0.5710 0.6790 2.4610 2.6650 ;
    LAYER PO ;
      RECT 2.9490 0.1030 2.9790 1.6210 ;
      RECT 2.7970 0.1030 2.8270 1.6210 ;
      RECT 2.6450 0.1030 2.6750 1.6210 ;
      RECT 2.4930 0.1030 2.5230 1.6210 ;
      RECT 0.0610 0.1030 0.0910 1.6210 ;
      RECT 0.2130 0.1030 0.2430 1.6210 ;
      RECT 0.3650 0.1030 0.3950 1.6210 ;
      RECT 0.5170 0.1030 0.5470 1.6210 ;
      RECT 0.5170 1.7330 0.5470 3.2510 ;
      RECT 0.3650 1.7330 0.3950 3.2510 ;
      RECT 0.2130 1.7330 0.2430 3.2510 ;
      RECT 0.0610 1.7330 0.0910 3.2510 ;
      RECT 2.4930 1.7330 2.5230 3.2510 ;
      RECT 2.6450 1.7330 2.6750 3.2510 ;
      RECT 2.7970 1.7330 2.8270 3.2510 ;
      RECT 2.9490 1.7330 2.9790 3.2510 ;
      RECT 1.2770 1.7330 1.3070 3.2510 ;
      RECT 1.1250 1.7330 1.1550 3.2510 ;
      RECT 1.7330 1.7330 1.7630 3.2510 ;
      RECT 1.4290 1.7330 1.4590 3.2510 ;
      RECT 0.9730 1.7330 1.0030 3.2510 ;
      RECT 0.8210 1.7330 0.8510 3.2510 ;
      RECT 1.5810 1.7330 1.6110 3.2510 ;
      RECT 0.6690 1.7330 0.6990 3.2510 ;
      RECT 1.8850 1.7330 1.9150 3.2510 ;
      RECT 2.0370 1.7330 2.0670 3.2510 ;
      RECT 2.1890 1.7330 2.2190 3.2510 ;
      RECT 2.3410 1.7330 2.3710 3.2510 ;
      RECT 2.3410 0.1030 2.3710 1.6210 ;
      RECT 2.1890 0.1030 2.2190 1.6210 ;
      RECT 2.0370 0.1030 2.0670 1.6210 ;
      RECT 1.8850 0.1030 1.9150 1.6210 ;
      RECT 0.6690 0.1030 0.6990 1.6210 ;
      RECT 1.5810 0.1030 1.6110 1.6210 ;
      RECT 0.8210 0.1030 0.8510 1.6210 ;
      RECT 0.9730 0.1030 1.0030 1.6210 ;
      RECT 1.4290 0.1030 1.4590 1.6210 ;
      RECT 1.7330 0.1030 1.7630 1.6210 ;
      RECT 1.1250 0.1030 1.1550 1.6210 ;
      RECT 1.2770 0.1030 1.3070 1.6210 ;
  END
END HEADX8_LVT

MACRO IBUFFX16_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.952 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.9520 1.7020 ;
        RECT 0.4310 0.9920 0.4810 1.6420 ;
        RECT 0.7350 0.9920 0.7850 1.6420 ;
        RECT 3.4710 0.9920 3.5210 1.6420 ;
        RECT 1.0390 0.9920 1.0890 1.6420 ;
        RECT 3.1670 0.9920 3.2170 1.6420 ;
        RECT 2.8630 0.9920 2.9130 1.6420 ;
        RECT 2.5590 0.9920 2.6090 1.6420 ;
        RECT 1.9510 0.9920 2.0010 1.6420 ;
        RECT 2.2550 0.9920 2.3050 1.6420 ;
        RECT 1.6470 0.9920 1.6970 1.6420 ;
        RECT 1.3430 0.9920 1.3930 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.9520 0.0300 ;
        RECT 0.4310 0.0300 0.4810 0.4100 ;
        RECT 0.7350 0.0300 0.7850 0.4100 ;
        RECT 3.4710 0.0300 3.5210 0.4100 ;
        RECT 3.1670 0.0300 3.2170 0.4100 ;
        RECT 1.0390 0.0300 1.0890 0.4100 ;
        RECT 2.8630 0.0300 2.9130 0.4100 ;
        RECT 2.5590 0.0300 2.6090 0.4100 ;
        RECT 1.9510 0.0300 2.0010 0.4100 ;
        RECT 2.2550 0.0300 2.3050 0.4100 ;
        RECT 1.6470 0.0300 1.6970 0.4100 ;
        RECT 1.3430 0.0300 1.3930 0.4100 ;
    END
  END VSS

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6600 0.4360 0.7100 ;
        RECT 0.2490 0.7100 0.3620 0.8150 ;
    END
    ANTENNAGATEAREA 0.0366 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1910 0.5370 3.8550 0.5870 ;
        RECT 3.6820 0.5870 3.8550 0.6630 ;
        RECT 3.6230 0.1160 3.6730 0.5370 ;
        RECT 3.3190 0.1160 3.3690 0.5370 ;
        RECT 2.1030 0.1160 2.1530 0.5370 ;
        RECT 2.4070 0.1170 2.4570 0.5370 ;
        RECT 2.7110 0.1160 2.7610 0.5370 ;
        RECT 3.0150 0.1160 3.0650 0.5370 ;
        RECT 1.7990 0.1160 1.8490 0.5370 ;
        RECT 1.1910 0.1160 1.2410 0.5370 ;
        RECT 1.4950 0.1160 1.5450 0.5370 ;
        RECT 3.6820 0.6630 3.7320 0.8920 ;
        RECT 1.1910 0.8920 3.7320 0.9420 ;
        RECT 3.6230 0.9420 3.6730 1.5640 ;
        RECT 3.3190 0.9420 3.3690 1.5640 ;
        RECT 3.0150 0.9420 3.0650 1.5640 ;
        RECT 2.1030 0.9420 2.1530 1.5640 ;
        RECT 2.4070 0.9420 2.4570 1.5650 ;
        RECT 2.7110 0.9420 2.7610 1.5640 ;
        RECT 1.1910 0.9420 1.2410 1.5640 ;
        RECT 1.4950 0.9420 1.5450 1.5640 ;
        RECT 1.7990 0.9420 1.8490 1.5640 ;
    END
    ANTENNADIFFAREA 1.2904 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 4.0670 1.7730 ;
    LAYER M1 ;
      RECT 1.0940 0.6600 3.6280 0.7100 ;
      RECT 0.5830 0.1160 0.6330 0.5370 ;
      RECT 0.5830 0.9420 0.6330 1.5640 ;
      RECT 0.8870 0.1160 0.9370 0.5370 ;
      RECT 0.8870 0.9420 0.9370 1.5640 ;
      RECT 1.0900 0.8740 1.1400 0.8920 ;
      RECT 0.5830 0.8920 1.1400 0.9420 ;
      RECT 1.0900 0.8420 1.1410 0.8740 ;
      RECT 1.0940 0.7100 1.1440 0.8420 ;
      RECT 1.0940 0.6370 1.1440 0.6600 ;
      RECT 1.0940 0.6330 1.1410 0.6370 ;
      RECT 0.5830 0.5370 1.1410 0.5870 ;
      RECT 1.0910 0.5870 1.1410 0.6330 ;
      RECT 0.4870 0.6600 1.0440 0.7100 ;
      RECT 0.2790 0.9420 0.3290 1.5640 ;
      RECT 0.2790 0.1160 0.3290 0.5370 ;
      RECT 0.4870 0.7100 0.5370 0.8320 ;
      RECT 0.4870 0.6420 0.5370 0.6600 ;
      RECT 0.4830 0.8320 0.5370 0.8700 ;
      RECT 0.4830 0.8700 0.5330 0.8920 ;
      RECT 0.4830 0.5870 0.5330 0.6070 ;
      RECT 0.2790 0.5370 0.5330 0.5870 ;
      RECT 0.2790 0.8920 0.5330 0.9420 ;
      RECT 0.4830 0.6070 0.5370 0.6100 ;
      RECT 0.4860 0.6100 0.5370 0.6420 ;
    LAYER PO ;
      RECT 3.8610 0.0690 3.8910 1.6060 ;
      RECT 3.5570 0.0690 3.5870 1.6060 ;
      RECT 2.3410 0.0690 2.3710 1.6060 ;
      RECT 2.4930 0.0690 2.5230 1.6060 ;
      RECT 2.6450 0.0690 2.6750 1.6060 ;
      RECT 3.2530 0.0690 3.2830 1.6060 ;
      RECT 3.1010 0.0690 3.1310 1.6060 ;
      RECT 2.9490 0.0690 2.9790 1.6060 ;
      RECT 2.7970 0.0690 2.8270 1.6060 ;
      RECT 3.4050 0.0690 3.4350 1.6060 ;
      RECT 2.1890 0.0690 2.2190 1.6060 ;
      RECT 2.0370 0.0690 2.0670 1.6060 ;
      RECT 1.8850 0.0690 1.9150 1.6060 ;
      RECT 1.1250 0.0690 1.1550 1.6060 ;
      RECT 1.2770 0.0690 1.3070 1.6060 ;
      RECT 1.7330 0.0690 1.7630 1.6060 ;
      RECT 1.5810 0.0690 1.6110 1.6060 ;
      RECT 1.4290 0.0690 1.4590 1.6060 ;
      RECT 0.0610 0.0710 0.0910 1.6060 ;
      RECT 0.8210 0.0690 0.8510 1.6060 ;
      RECT 0.9730 0.0690 1.0030 1.6060 ;
      RECT 0.3650 0.0690 0.3950 1.6060 ;
      RECT 0.6690 0.0690 0.6990 1.6060 ;
      RECT 0.2130 0.0710 0.2430 1.6060 ;
      RECT 0.5170 0.0710 0.5470 1.6060 ;
      RECT 3.7090 0.0690 3.7390 1.6060 ;
  END
END IBUFFX16_LVT

MACRO IBUFFX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.52 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6600 0.4360 0.7100 ;
        RECT 0.2490 0.7100 0.3620 0.8150 ;
    END
    ANTENNAGATEAREA 0.0186 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.5200 1.7020 ;
        RECT 0.2790 0.8650 0.3290 1.6420 ;
        RECT 0.5830 0.8930 0.6330 1.6420 ;
        RECT 1.0390 0.9920 1.0890 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.5200 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.5600 ;
        RECT 0.5830 0.0300 0.6330 0.5540 ;
        RECT 1.0390 0.0300 1.0890 0.4100 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8870 0.1160 0.9370 0.5370 ;
        RECT 0.8870 0.5370 1.4230 0.5870 ;
        RECT 1.2470 0.5870 1.4230 0.6630 ;
        RECT 1.1910 0.1160 1.2410 0.5370 ;
        RECT 1.2470 0.6630 1.2970 0.8920 ;
        RECT 0.8870 0.8920 1.2970 0.9420 ;
        RECT 1.1910 0.9420 1.2410 1.5640 ;
        RECT 0.8870 0.9420 0.9370 1.5640 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.6350 1.7730 ;
    LAYER M1 ;
      RECT 0.4870 0.6600 0.7400 0.7100 ;
      RECT 0.4870 0.7100 0.5370 0.7750 ;
      RECT 0.4870 0.6300 0.5370 0.6600 ;
      RECT 0.4310 0.7750 0.5370 0.8250 ;
      RECT 0.4830 0.6070 0.5370 0.6100 ;
      RECT 0.4860 0.6100 0.5370 0.6300 ;
      RECT 0.4830 0.5820 0.5330 0.6070 ;
      RECT 0.4310 0.5320 0.5330 0.5820 ;
      RECT 0.4310 0.8250 0.4810 1.1650 ;
      RECT 0.4310 0.3620 0.4810 0.5320 ;
      RECT 0.7910 0.6600 1.1960 0.7100 ;
      RECT 0.7350 0.8260 0.7850 1.1910 ;
      RECT 0.7350 0.2850 0.7850 0.5320 ;
      RECT 0.7910 0.7100 0.8410 0.7760 ;
      RECT 0.7910 0.6410 0.8410 0.6600 ;
      RECT 0.7350 0.7760 0.8410 0.8260 ;
      RECT 0.7870 0.6370 0.8410 0.6410 ;
      RECT 0.7350 0.5320 0.8370 0.5820 ;
      RECT 0.7870 0.5820 0.8370 0.6370 ;
    LAYER PO ;
      RECT 0.0610 0.0690 0.0910 1.6060 ;
      RECT 0.2130 0.0690 0.2430 1.6060 ;
      RECT 0.3650 0.0710 0.3950 1.6060 ;
      RECT 0.6690 0.0690 0.6990 1.6060 ;
      RECT 0.5170 0.0710 0.5470 1.6060 ;
      RECT 0.8210 0.0710 0.8510 1.6060 ;
      RECT 0.9730 0.0690 1.0030 1.6060 ;
      RECT 1.4290 0.0710 1.4590 1.6060 ;
      RECT 1.2770 0.0710 1.3070 1.6060 ;
      RECT 1.1250 0.0690 1.1550 1.6060 ;
  END
END IBUFFX2_LVT

MACRO IBUFFX32_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.992 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6600 0.5880 0.7100 ;
        RECT 0.2490 0.7100 0.3620 0.8150 ;
    END
    ANTENNAGATEAREA 0.0732 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 6.9920 1.7020 ;
        RECT 2.5590 0.9920 2.6090 1.6420 ;
        RECT 2.8630 0.9920 2.9130 1.6420 ;
        RECT 2.2550 0.9920 2.3050 1.6420 ;
        RECT 1.9510 0.9920 2.0010 1.6420 ;
        RECT 1.0390 0.9920 1.0890 1.6420 ;
        RECT 0.4310 0.9920 0.4810 1.6420 ;
        RECT 1.3430 0.9920 1.3930 1.6420 ;
        RECT 1.6470 0.9920 1.6970 1.6420 ;
        RECT 6.5110 0.9920 6.5610 1.6420 ;
        RECT 6.2070 0.9920 6.2570 1.6420 ;
        RECT 5.9030 0.9920 5.9530 1.6420 ;
        RECT 5.5990 0.9920 5.6490 1.6420 ;
        RECT 5.2950 0.9920 5.3450 1.6420 ;
        RECT 4.9910 0.9920 5.0410 1.6420 ;
        RECT 4.6870 0.9920 4.7370 1.6420 ;
        RECT 4.3830 0.9920 4.4330 1.6420 ;
        RECT 4.0790 0.9920 4.1290 1.6420 ;
        RECT 3.7750 0.9920 3.8250 1.6420 ;
        RECT 0.7350 0.9920 0.7850 1.6420 ;
        RECT 3.4710 0.9920 3.5210 1.6420 ;
        RECT 3.1670 0.9920 3.2170 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 6.9920 0.0300 ;
        RECT 2.5590 0.0300 2.6090 0.4100 ;
        RECT 2.8630 0.0300 2.9130 0.4100 ;
        RECT 2.2550 0.0300 2.3050 0.4100 ;
        RECT 1.9510 0.0300 2.0010 0.4100 ;
        RECT 0.4310 0.0300 0.4810 0.4100 ;
        RECT 1.0390 0.0300 1.0890 0.4100 ;
        RECT 1.3430 0.0300 1.3930 0.4100 ;
        RECT 1.6470 0.0300 1.6970 0.4100 ;
        RECT 6.5110 0.0300 6.5610 0.4100 ;
        RECT 6.2070 0.0300 6.2570 0.4100 ;
        RECT 5.9030 0.0300 5.9530 0.4100 ;
        RECT 5.5990 0.0300 5.6490 0.4100 ;
        RECT 5.2950 0.0300 5.3450 0.4100 ;
        RECT 4.9910 0.0300 5.0410 0.4100 ;
        RECT 4.6870 0.0300 4.7370 0.4100 ;
        RECT 4.3830 0.0300 4.4330 0.4100 ;
        RECT 0.7350 0.0300 0.7850 0.4100 ;
        RECT 4.0790 0.0300 4.1290 0.4100 ;
        RECT 3.7750 0.0300 3.8250 0.4100 ;
        RECT 3.4710 0.0300 3.5210 0.4100 ;
        RECT 3.1670 0.0300 3.2170 0.4100 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.5350 0.9420 4.5850 1.5640 ;
        RECT 4.8390 0.9420 4.8890 1.5640 ;
        RECT 5.1430 0.9420 5.1930 1.5640 ;
        RECT 5.4470 0.9420 5.4970 1.5640 ;
        RECT 5.7510 0.9420 5.8010 1.5640 ;
        RECT 6.0550 0.9420 6.1050 1.5640 ;
        RECT 6.3590 0.9420 6.4090 1.5640 ;
        RECT 6.6630 0.9420 6.7130 1.5640 ;
        RECT 3.0150 0.9420 3.0650 1.5650 ;
        RECT 3.6230 0.9420 3.6730 1.5640 ;
        RECT 3.9270 0.9420 3.9770 1.5640 ;
        RECT 4.2310 0.9420 4.2810 1.5640 ;
        RECT 2.4070 0.9420 2.4570 1.5640 ;
        RECT 2.1030 0.9420 2.1530 1.5640 ;
        RECT 1.7990 0.9420 1.8490 1.5640 ;
        RECT 3.3190 0.9420 3.3690 1.5640 ;
        RECT 2.7110 0.9420 2.7610 1.5640 ;
        RECT 1.7990 0.8920 6.7720 0.9420 ;
        RECT 6.7220 0.6630 6.7720 0.8920 ;
        RECT 1.7990 0.5370 6.8950 0.5870 ;
        RECT 2.7110 0.1160 2.7610 0.5370 ;
        RECT 3.9270 0.1160 3.9770 0.5370 ;
        RECT 4.2310 0.1160 4.2810 0.5370 ;
        RECT 2.1030 0.1160 2.1530 0.5370 ;
        RECT 1.7990 0.1160 1.8490 0.5370 ;
        RECT 2.4070 0.1160 2.4570 0.5370 ;
        RECT 3.6230 0.1160 3.6730 0.5370 ;
        RECT 3.3190 0.1160 3.3690 0.5370 ;
        RECT 3.0150 0.1170 3.0650 0.5370 ;
        RECT 6.7220 0.5870 6.8950 0.6630 ;
        RECT 4.5350 0.1160 4.5850 0.5370 ;
        RECT 4.8390 0.1160 4.8890 0.5370 ;
        RECT 5.1430 0.1160 5.1930 0.5370 ;
        RECT 5.4470 0.1160 5.4970 0.5370 ;
        RECT 5.7510 0.1160 5.8010 0.5370 ;
        RECT 6.0550 0.1160 6.1050 0.5370 ;
        RECT 6.3590 0.1160 6.4090 0.5370 ;
        RECT 6.6630 0.1160 6.7130 0.5370 ;
    END
    ANTENNADIFFAREA 2.4808 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 7.1070 1.7730 ;
    LAYER M1 ;
      RECT 1.7020 0.6600 6.6680 0.7100 ;
      RECT 0.8870 0.9420 0.9370 1.5640 ;
      RECT 0.8870 0.1160 0.9370 0.5370 ;
      RECT 1.1910 0.9420 1.2410 1.5640 ;
      RECT 1.1910 0.1160 1.2410 0.5370 ;
      RECT 1.4950 0.9420 1.5450 1.5640 ;
      RECT 1.4950 0.1160 1.5450 0.5370 ;
      RECT 1.7020 0.7100 1.7520 0.8180 ;
      RECT 1.6990 0.8180 1.7520 0.8420 ;
      RECT 0.8870 0.8920 1.7490 0.9420 ;
      RECT 1.6990 0.8420 1.7490 0.8920 ;
      RECT 1.7020 0.6370 1.7520 0.6600 ;
      RECT 1.7020 0.6310 1.7490 0.6370 ;
      RECT 0.8870 0.5370 1.7490 0.5870 ;
      RECT 1.6990 0.5870 1.7490 0.6310 ;
      RECT 0.6390 0.6600 1.6520 0.7100 ;
      RECT 0.2790 0.1160 0.3290 0.5370 ;
      RECT 0.2790 0.9420 0.3290 1.5640 ;
      RECT 0.5830 0.1160 0.6330 0.5370 ;
      RECT 0.5830 0.9420 0.6330 1.5640 ;
      RECT 0.6390 0.5870 0.6890 0.6600 ;
      RECT 0.6390 0.7100 0.6890 0.8920 ;
      RECT 0.2790 0.5370 0.6890 0.5870 ;
      RECT 0.2790 0.8920 0.6890 0.9420 ;
    LAYER PO ;
      RECT 6.4450 0.0690 6.4750 1.6060 ;
      RECT 6.1410 0.0690 6.1710 1.6060 ;
      RECT 6.2930 0.0690 6.3230 1.6060 ;
      RECT 5.8370 0.0690 5.8670 1.6060 ;
      RECT 5.9890 0.0690 6.0190 1.6060 ;
      RECT 5.6850 0.0690 5.7150 1.6060 ;
      RECT 5.5330 0.0690 5.5630 1.6060 ;
      RECT 5.3810 0.0690 5.4110 1.6060 ;
      RECT 5.2290 0.0690 5.2590 1.6060 ;
      RECT 4.9250 0.0690 4.9550 1.6060 ;
      RECT 5.0770 0.0690 5.1070 1.6060 ;
      RECT 4.3170 0.0690 4.3470 1.6060 ;
      RECT 4.4690 0.0690 4.4990 1.6060 ;
      RECT 4.1650 0.0690 4.1950 1.6060 ;
      RECT 4.6210 0.0690 4.6510 1.6060 ;
      RECT 4.7730 0.0690 4.8030 1.6060 ;
      RECT 2.9490 0.0690 2.9790 1.6060 ;
      RECT 3.1010 0.0690 3.1310 1.6060 ;
      RECT 3.2530 0.0690 3.2830 1.6060 ;
      RECT 3.8610 0.0690 3.8910 1.6060 ;
      RECT 3.7090 0.0690 3.7390 1.6060 ;
      RECT 3.5570 0.0690 3.5870 1.6060 ;
      RECT 3.4050 0.0690 3.4350 1.6060 ;
      RECT 4.0130 0.0690 4.0430 1.6060 ;
      RECT 2.7970 0.0690 2.8270 1.6060 ;
      RECT 2.6450 0.0690 2.6750 1.6060 ;
      RECT 2.4930 0.0690 2.5230 1.6060 ;
      RECT 1.7330 0.0690 1.7630 1.6060 ;
      RECT 1.8850 0.0690 1.9150 1.6060 ;
      RECT 2.3410 0.0690 2.3710 1.6060 ;
      RECT 2.1890 0.0690 2.2190 1.6060 ;
      RECT 2.0370 0.0690 2.0670 1.6060 ;
      RECT 0.0610 0.0710 0.0910 1.6060 ;
      RECT 0.6690 0.0690 0.6990 1.6060 ;
      RECT 0.5170 0.0690 0.5470 1.6060 ;
      RECT 1.1250 0.0690 1.1550 1.6060 ;
      RECT 1.2770 0.0690 1.3070 1.6060 ;
      RECT 1.4290 0.0690 1.4590 1.6060 ;
      RECT 0.9730 0.0690 1.0030 1.6060 ;
      RECT 0.8210 0.0690 0.8510 1.6060 ;
      RECT 1.5810 0.0690 1.6110 1.6060 ;
      RECT 0.2130 0.0710 0.2430 1.6060 ;
      RECT 0.3650 0.0690 0.3950 1.6060 ;
      RECT 6.9010 0.0690 6.9310 1.6060 ;
      RECT 6.7490 0.0690 6.7790 1.6060 ;
      RECT 6.5970 0.0690 6.6270 1.6060 ;
  END
END IBUFFX32_LVT

MACRO IBUFFX4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.824 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6600 0.4360 0.7100 ;
        RECT 0.2490 0.7100 0.3620 0.8150 ;
    END
    ANTENNAGATEAREA 0.0186 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.8240 1.7020 ;
        RECT 0.2790 0.8650 0.3290 1.6420 ;
        RECT 0.5830 0.9870 0.6330 1.6420 ;
        RECT 1.3430 0.9920 1.3930 1.6420 ;
        RECT 1.0390 0.9920 1.0890 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.8240 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.5590 ;
        RECT 0.5830 0.0300 0.6330 0.4050 ;
        RECT 1.3430 0.0300 1.3930 0.4100 ;
        RECT 1.0390 0.0300 1.0890 0.4100 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8870 0.5370 1.7270 0.5870 ;
        RECT 1.5500 0.5870 1.7270 0.6630 ;
        RECT 1.4950 0.1160 1.5450 0.5370 ;
        RECT 0.8870 0.1160 0.9370 0.5370 ;
        RECT 1.1910 0.1160 1.2410 0.5370 ;
        RECT 1.5500 0.6630 1.6000 0.8920 ;
        RECT 0.8870 0.8920 1.6000 0.9420 ;
        RECT 0.8870 0.9420 0.9370 1.5640 ;
        RECT 1.1910 0.9420 1.2410 1.5640 ;
        RECT 1.4950 0.9420 1.5450 1.5640 ;
    END
    ANTENNADIFFAREA 0.3976 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1120 0.6790 1.9390 1.7730 ;
    LAYER M1 ;
      RECT 0.4870 0.6600 0.7400 0.7100 ;
      RECT 0.4870 0.6370 0.5370 0.6600 ;
      RECT 0.4870 0.7100 0.5370 0.8220 ;
      RECT 0.4310 0.8220 0.5370 0.8720 ;
      RECT 0.4830 0.5820 0.5330 0.6090 ;
      RECT 0.4310 0.5320 0.5330 0.5820 ;
      RECT 0.4830 0.6090 0.5370 0.6100 ;
      RECT 0.4860 0.6100 0.5370 0.6370 ;
      RECT 0.4310 0.8720 0.4810 1.1180 ;
      RECT 0.4310 0.3540 0.4810 0.5320 ;
      RECT 0.7910 0.6600 1.5000 0.7100 ;
      RECT 0.7350 0.8720 0.7850 1.5590 ;
      RECT 0.7350 0.1110 0.7850 0.5320 ;
      RECT 0.7910 0.7100 0.8410 0.8220 ;
      RECT 0.7350 0.8220 0.8410 0.8420 ;
      RECT 0.7350 0.8420 0.8370 0.8720 ;
      RECT 0.7910 0.6370 0.8410 0.6600 ;
      RECT 0.7350 0.5320 0.8370 0.5820 ;
      RECT 0.7870 0.5820 0.8370 0.6370 ;
    LAYER PO ;
      RECT 0.3650 0.0690 0.3950 1.6060 ;
      RECT 0.0610 0.0710 0.0910 1.6060 ;
      RECT 0.6690 0.0690 0.6990 1.6060 ;
      RECT 0.2130 0.0710 0.2430 1.6060 ;
      RECT 0.5170 0.0710 0.5470 1.6060 ;
      RECT 1.7330 0.0650 1.7630 1.6000 ;
      RECT 1.5810 0.0650 1.6110 1.6000 ;
      RECT 0.8210 0.0710 0.8510 1.6060 ;
      RECT 0.9730 0.0690 1.0030 1.6060 ;
      RECT 1.4290 0.0690 1.4590 1.6060 ;
      RECT 1.2770 0.0690 1.3070 1.6060 ;
      RECT 1.1250 0.0690 1.1550 1.6060 ;
  END
END IBUFFX4_LVT

MACRO IBUFFX8_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.584 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6800 0.4360 0.7300 ;
        RECT 0.2490 0.7300 0.3620 0.8150 ;
    END
    ANTENNAGATEAREA 0.0237 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.5840 1.7020 ;
        RECT 0.4310 0.9920 0.4810 1.6420 ;
        RECT 0.7350 0.9920 0.7850 1.6420 ;
        RECT 1.7990 0.9920 1.8490 1.6420 ;
        RECT 2.1030 0.9920 2.1530 1.6420 ;
        RECT 1.4950 0.9920 1.5450 1.6420 ;
        RECT 1.1910 0.9920 1.2410 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.5840 0.0300 ;
        RECT 0.4310 0.0300 0.4810 0.4870 ;
        RECT 0.7350 0.0300 0.7850 0.4100 ;
        RECT 1.7990 0.0300 1.8490 0.4100 ;
        RECT 2.1030 0.0300 2.1530 0.4100 ;
        RECT 1.4950 0.0300 1.5450 0.4100 ;
        RECT 1.1910 0.0300 1.2410 0.4100 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0390 0.5370 2.4870 0.5870 ;
        RECT 2.3110 0.5870 2.4870 0.6630 ;
        RECT 1.9510 0.1160 2.0010 0.5370 ;
        RECT 2.2550 0.1170 2.3050 0.5370 ;
        RECT 1.6470 0.1160 1.6970 0.5370 ;
        RECT 1.0390 0.1160 1.0890 0.5370 ;
        RECT 1.3430 0.1160 1.3930 0.5370 ;
        RECT 2.3110 0.6630 2.3610 0.8920 ;
        RECT 1.0390 0.8920 2.3610 0.9420 ;
        RECT 1.9510 0.9420 2.0010 1.5640 ;
        RECT 2.2550 0.9420 2.3050 1.5650 ;
        RECT 1.0390 0.9420 1.0890 1.5640 ;
        RECT 1.3430 0.9420 1.3930 1.5640 ;
        RECT 1.6470 0.9420 1.6970 1.5640 ;
    END
    ANTENNADIFFAREA 0.6952 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 2.6990 1.7730 ;
    LAYER M1 ;
      RECT 0.9430 0.6600 2.2600 0.7100 ;
      RECT 0.5830 0.9420 0.6330 1.5640 ;
      RECT 0.5830 0.1160 0.6330 0.5370 ;
      RECT 0.8870 0.9420 0.9370 1.5640 ;
      RECT 0.8870 0.1160 0.9370 0.5370 ;
      RECT 0.9430 0.6420 0.9930 0.6600 ;
      RECT 0.9430 0.7100 0.9930 0.8420 ;
      RECT 0.9430 0.8420 0.9890 0.8500 ;
      RECT 0.5830 0.8920 0.9890 0.9420 ;
      RECT 0.9390 0.8500 0.9890 0.8920 ;
      RECT 0.9390 0.6370 0.9930 0.6420 ;
      RECT 0.5830 0.5370 0.9890 0.5870 ;
      RECT 0.9390 0.5870 0.9890 0.6370 ;
      RECT 0.4870 0.6600 0.8920 0.7100 ;
      RECT 0.2790 0.3050 0.3290 0.5370 ;
      RECT 0.2790 0.9420 0.3290 1.2880 ;
      RECT 0.4870 0.6490 0.5370 0.6600 ;
      RECT 0.4870 0.7100 0.5370 0.8110 ;
      RECT 0.4830 0.8110 0.5370 0.8700 ;
      RECT 0.4830 0.5870 0.5330 0.6090 ;
      RECT 0.4830 0.8700 0.5330 0.8920 ;
      RECT 0.4830 0.6090 0.5370 0.6300 ;
      RECT 0.4860 0.6300 0.5370 0.6490 ;
      RECT 0.2790 0.8920 0.5330 0.9420 ;
      RECT 0.2790 0.5370 0.5330 0.5870 ;
    LAYER PO ;
      RECT 0.0610 0.0710 0.0910 1.6060 ;
      RECT 0.3650 0.0690 0.3950 1.6060 ;
      RECT 0.2130 0.0710 0.2430 1.6060 ;
      RECT 0.8210 0.0690 0.8510 1.6060 ;
      RECT 2.1890 0.0690 2.2190 1.6060 ;
      RECT 2.3410 0.0690 2.3710 1.6060 ;
      RECT 2.4930 0.0690 2.5230 1.6060 ;
      RECT 0.5170 0.0710 0.5470 1.6060 ;
      RECT 0.6690 0.0690 0.6990 1.6060 ;
      RECT 2.0370 0.0690 2.0670 1.6060 ;
      RECT 1.8850 0.0690 1.9150 1.6060 ;
      RECT 1.7330 0.0690 1.7630 1.6060 ;
      RECT 0.9730 0.0690 1.0030 1.6060 ;
      RECT 1.1250 0.0690 1.1550 1.6060 ;
      RECT 1.5810 0.0690 1.6110 1.6060 ;
      RECT 1.4290 0.0690 1.4590 1.6060 ;
      RECT 1.2770 0.0690 1.3070 1.6060 ;
  END
END IBUFFX8_LVT

MACRO INVX0_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.76 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6800 0.4210 0.7300 ;
        RECT 0.2490 0.7300 0.3620 0.8150 ;
    END
    ANTENNAGATEAREA 0.0237 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 0.7600 1.7020 ;
        RECT 0.2790 0.9280 0.3290 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 0.7600 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.5640 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4310 0.3050 0.4810 0.5370 ;
        RECT 0.4310 0.5370 0.6630 0.5870 ;
        RECT 0.4710 0.5870 0.6630 0.6630 ;
        RECT 0.4710 0.6630 0.5210 0.8230 ;
        RECT 0.4310 0.8230 0.5210 0.8730 ;
        RECT 0.4310 0.8730 0.4810 1.2880 ;
    END
    ANTENNADIFFAREA 0.0805 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 0.8750 1.7730 ;
    LAYER PO ;
      RECT 0.2130 0.0710 0.2430 1.6060 ;
      RECT 0.3650 0.0690 0.3950 1.6060 ;
      RECT 0.6690 0.0710 0.6990 1.6060 ;
      RECT 0.5170 0.0710 0.5470 1.6060 ;
      RECT 0.0610 0.0710 0.0910 1.6060 ;
  END
END INVX0_LVT

MACRO INVX16_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.04 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6600 2.7160 0.7100 ;
        RECT 0.2490 0.7100 0.3620 0.8150 ;
    END
    ANTENNAGATEAREA 0.5856 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.0400 1.7020 ;
        RECT 2.5590 0.9920 2.6090 1.6420 ;
        RECT 2.2550 0.9920 2.3050 1.6420 ;
        RECT 1.9510 0.9920 2.0010 1.6420 ;
        RECT 1.6470 0.9920 1.6970 1.6420 ;
        RECT 1.0390 0.9920 1.0890 1.6420 ;
        RECT 1.3430 0.9920 1.3930 1.6420 ;
        RECT 0.7350 0.9920 0.7850 1.6420 ;
        RECT 0.4310 0.9920 0.4810 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.0400 0.0300 ;
        RECT 2.5590 0.0300 2.6090 0.4100 ;
        RECT 2.2550 0.0300 2.3050 0.4100 ;
        RECT 1.9510 0.0300 2.0010 0.4100 ;
        RECT 1.6470 0.0300 1.6970 0.4100 ;
        RECT 1.0390 0.0300 1.0890 0.4100 ;
        RECT 1.3430 0.0300 1.3930 0.4100 ;
        RECT 0.7350 0.0300 0.7850 0.4100 ;
        RECT 0.4310 0.0300 0.4810 0.4100 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2790 0.5370 2.9430 0.5870 ;
        RECT 2.7700 0.5870 2.9430 0.6630 ;
        RECT 2.7110 0.1160 2.7610 0.5370 ;
        RECT 2.4070 0.1160 2.4570 0.5370 ;
        RECT 1.1910 0.1160 1.2410 0.5370 ;
        RECT 1.4950 0.1170 1.5450 0.5370 ;
        RECT 1.7990 0.1160 1.8490 0.5370 ;
        RECT 2.1030 0.1160 2.1530 0.5370 ;
        RECT 0.8870 0.1160 0.9370 0.5370 ;
        RECT 0.2790 0.1160 0.3290 0.5370 ;
        RECT 0.5830 0.1160 0.6330 0.5370 ;
        RECT 2.7700 0.6630 2.8200 0.8920 ;
        RECT 0.2790 0.8920 2.8200 0.9420 ;
        RECT 2.7110 0.9420 2.7610 1.5640 ;
        RECT 2.4070 0.9420 2.4570 1.5640 ;
        RECT 2.1030 0.9420 2.1530 1.5640 ;
        RECT 1.1910 0.9420 1.2410 1.5640 ;
        RECT 1.4950 0.9420 1.5450 1.5650 ;
        RECT 1.7990 0.9420 1.8490 1.5640 ;
        RECT 0.2790 0.9420 0.3290 1.5640 ;
        RECT 0.5830 0.9420 0.6330 1.5640 ;
        RECT 0.8870 0.9420 0.9370 1.5640 ;
    END
    ANTENNADIFFAREA 1.2904 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 3.1550 1.7730 ;
    LAYER PO ;
      RECT 2.7970 0.0690 2.8270 1.6060 ;
      RECT 2.9490 0.0690 2.9790 1.6060 ;
      RECT 2.6450 0.0690 2.6750 1.6060 ;
      RECT 1.4290 0.0690 1.4590 1.6060 ;
      RECT 1.5810 0.0690 1.6110 1.6060 ;
      RECT 1.7330 0.0690 1.7630 1.6060 ;
      RECT 2.3410 0.0690 2.3710 1.6060 ;
      RECT 2.1890 0.0690 2.2190 1.6060 ;
      RECT 2.0370 0.0690 2.0670 1.6060 ;
      RECT 1.8850 0.0690 1.9150 1.6060 ;
      RECT 2.4930 0.0690 2.5230 1.6060 ;
      RECT 1.2770 0.0690 1.3070 1.6060 ;
      RECT 1.1250 0.0690 1.1550 1.6060 ;
      RECT 0.9730 0.0690 1.0030 1.6060 ;
      RECT 0.2130 0.0690 0.2430 1.6060 ;
      RECT 0.3650 0.0690 0.3950 1.6060 ;
      RECT 0.8210 0.0690 0.8510 1.6060 ;
      RECT 0.6690 0.0690 0.6990 1.6060 ;
      RECT 0.5170 0.0690 0.5470 1.6060 ;
      RECT 0.0610 0.0690 0.0910 1.6060 ;
  END
END INVX16_LVT

MACRO INVX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.76 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6600 0.4210 0.7100 ;
        RECT 0.2490 0.7100 0.3620 0.8150 ;
    END
    ANTENNAGATEAREA 0.0366 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 0.7600 1.7020 ;
        RECT 0.4310 0.9920 0.4810 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 0.7600 0.0300 ;
        RECT 0.4310 0.0300 0.4810 0.4100 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2790 0.1160 0.3290 0.5370 ;
        RECT 0.2790 0.5370 0.6630 0.5870 ;
        RECT 0.4710 0.5870 0.6630 0.6630 ;
        RECT 0.4710 0.6630 0.5210 0.8920 ;
        RECT 0.2790 0.8920 0.5210 0.9420 ;
        RECT 0.2790 0.9420 0.3290 1.5640 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 0.8750 1.7730 ;
    LAYER PO ;
      RECT 0.2130 0.0710 0.2430 1.6060 ;
      RECT 0.3650 0.0690 0.3950 1.6060 ;
      RECT 0.6690 0.0710 0.6990 1.6060 ;
      RECT 0.5170 0.0710 0.5470 1.6060 ;
      RECT 0.0610 0.0710 0.0910 1.6060 ;
  END
END INVX1_LVT

MACRO INVX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.912 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6600 0.5880 0.7100 ;
        RECT 0.2490 0.7100 0.3620 0.8150 ;
    END
    ANTENNAGATEAREA 0.0732 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 0.9120 1.7020 ;
        RECT 0.4310 0.9920 0.4810 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 0.9120 0.0300 ;
        RECT 0.4310 0.0300 0.4810 0.4100 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2790 0.1160 0.3290 0.5370 ;
        RECT 0.2790 0.5370 0.8150 0.5870 ;
        RECT 0.6390 0.5870 0.8150 0.6630 ;
        RECT 0.5830 0.1160 0.6330 0.5370 ;
        RECT 0.6390 0.6630 0.6890 0.8920 ;
        RECT 0.2790 0.8920 0.6890 0.9420 ;
        RECT 0.5830 0.9420 0.6330 1.5640 ;
        RECT 0.2790 0.9420 0.3290 1.5640 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.0270 1.7730 ;
    LAYER PO ;
      RECT 0.2130 0.0710 0.2430 1.6060 ;
      RECT 0.3650 0.0690 0.3950 1.6060 ;
      RECT 0.8210 0.0710 0.8510 1.6060 ;
      RECT 0.6690 0.0710 0.6990 1.6060 ;
      RECT 0.5170 0.0690 0.5470 1.6060 ;
      RECT 0.0610 0.0710 0.0910 1.6060 ;
  END
END INVX2_LVT

MACRO FOOTX16_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.256 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VSSG
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.6660 1.0090 0.8560 1.1190 ;
        RECT 0.7350 1.1190 0.7850 1.1650 ;
        RECT 0.7350 0.8810 0.7850 1.0090 ;
        RECT 0.7350 0.8310 3.3690 0.8810 ;
        RECT 1.4950 0.8810 1.5450 1.5610 ;
        RECT 3.3190 0.8810 3.3690 1.5610 ;
        RECT 1.1910 0.8810 1.2410 1.5610 ;
        RECT 2.1030 0.8810 2.1530 1.5610 ;
        RECT 2.4070 0.8810 2.4570 1.5610 ;
        RECT 2.7110 0.8810 2.7610 1.5610 ;
        RECT 3.0150 0.8810 3.0650 1.5610 ;
        RECT 1.7990 0.8810 1.8490 1.5610 ;
    END
  END VSSG

  PIN VSS
    DIRECTION OUTPUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.2560 1.7020 ;
        RECT 1.0390 1.2010 1.0890 1.6420 ;
        RECT 1.6470 1.2010 1.6970 1.6420 ;
        RECT 1.3430 1.2010 1.3930 1.6420 ;
        RECT 3.4710 1.2010 3.5210 1.6420 ;
        RECT 3.1670 1.2010 3.2170 1.6420 ;
        RECT 2.8630 1.2010 2.9130 1.6420 ;
        RECT 2.5590 1.2010 2.6090 1.6420 ;
        RECT 2.2550 1.2010 2.3050 1.6420 ;
        RECT 1.9510 1.2010 2.0010 1.6420 ;
    END
  END VSS

  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0990 0.6700 3.4610 0.7300 ;
        RECT 1.1200 0.5530 1.3100 0.6700 ;
    END
    ANTENNAGATEAREA 0.2016 ;
  END SLEEP

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.2560 0.0300 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 4.2560 3.3740 ;
    END
  END VDD
  OBS
    LAYER NWELL ;
      RECT -0.1120 2.3510 4.3850 3.4540 ;
      RECT 0.2300 1.6770 4.0260 2.3510 ;
      RECT 0.2300 0.9930 0.5620 1.6770 ;
      RECT 3.6620 0.9930 4.0260 1.6770 ;
      RECT -0.1090 0.7460 0.5620 0.9930 ;
      RECT 3.6620 0.7460 4.3830 0.9930 ;
      RECT -0.1090 -0.1410 4.3830 0.7460 ;
    LAYER PO ;
      RECT 1.8850 2.0450 1.9150 3.1790 ;
      RECT 2.1890 2.0450 2.2190 3.1790 ;
      RECT 1.2770 2.0450 1.3070 3.1790 ;
      RECT 2.3410 2.0450 2.3710 3.1790 ;
      RECT 1.1250 2.0450 1.1550 3.1790 ;
      RECT 1.7330 2.0450 1.7630 3.1790 ;
      RECT 1.4290 2.0450 1.4590 3.1790 ;
      RECT 0.9730 2.0450 1.0030 3.1790 ;
      RECT 3.7090 2.0450 3.7390 3.1790 ;
      RECT 0.8210 2.0450 0.8510 3.1790 ;
      RECT 1.5810 2.0450 1.6110 3.1790 ;
      RECT 0.6690 2.0450 0.6990 3.1790 ;
      RECT 2.0370 2.0450 2.0670 3.1790 ;
      RECT 3.5570 2.0450 3.5870 3.1790 ;
      RECT 3.4050 2.0450 3.4350 3.1790 ;
      RECT 3.2530 2.0450 3.2830 3.1790 ;
      RECT 3.1010 2.0450 3.1310 3.1790 ;
      RECT 2.9490 2.0450 2.9790 3.1790 ;
      RECT 2.7970 2.0450 2.8270 3.1790 ;
      RECT 2.6450 2.0450 2.6750 3.1790 ;
      RECT 2.4930 2.0450 2.5230 3.1790 ;
      RECT 4.1650 2.0450 4.1950 3.1790 ;
      RECT 4.0130 2.0450 4.0430 3.1790 ;
      RECT 3.8610 2.0450 3.8910 3.1790 ;
      RECT 0.3650 2.0450 0.3950 3.1790 ;
      RECT 0.2130 2.0450 0.2430 3.1790 ;
      RECT 0.0610 2.0450 0.0910 3.1790 ;
      RECT 0.5170 2.0450 0.5470 3.1790 ;
      RECT 0.6690 0.4870 0.6990 1.6210 ;
      RECT 0.5170 0.4870 0.5470 1.6210 ;
      RECT 0.3650 0.4870 0.3950 1.6210 ;
      RECT 0.0610 0.4870 0.0910 1.6210 ;
      RECT 0.2130 0.4870 0.2430 1.6210 ;
      RECT 4.0130 0.4870 4.0430 1.6210 ;
      RECT 3.8610 0.4870 3.8910 1.6210 ;
      RECT 4.1650 0.4870 4.1950 1.6210 ;
      RECT 2.4930 0.4870 2.5230 1.6210 ;
      RECT 2.6450 0.4870 2.6750 1.6210 ;
      RECT 2.7970 0.4870 2.8270 1.6210 ;
      RECT 2.9490 0.4870 2.9790 1.6210 ;
      RECT 3.1010 0.4870 3.1310 1.6210 ;
      RECT 3.2530 0.4870 3.2830 1.6210 ;
      RECT 3.4050 0.4870 3.4350 1.6210 ;
      RECT 3.5570 0.4870 3.5870 1.6210 ;
      RECT 2.0370 0.4870 2.0670 1.6210 ;
      RECT 1.5810 0.4870 1.6110 1.6210 ;
      RECT 0.8210 0.4870 0.8510 1.6210 ;
      RECT 3.7090 0.4870 3.7390 1.6210 ;
      RECT 0.9730 0.4870 1.0030 1.6210 ;
      RECT 1.4290 0.4870 1.4590 1.6210 ;
      RECT 1.7330 0.4870 1.7630 1.6210 ;
      RECT 1.1250 0.4870 1.1550 1.6210 ;
      RECT 2.3410 0.4870 2.3710 1.6210 ;
      RECT 1.2770 0.4870 1.3070 1.6210 ;
      RECT 2.1890 0.4870 2.2190 1.6210 ;
      RECT 1.8850 0.4870 1.9150 1.6210 ;
  END
END FOOTX16_LVT

MACRO FOOTX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.128 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VSSG
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.6660 1.0090 0.8560 1.1190 ;
        RECT 0.7350 1.1190 0.7850 1.1650 ;
        RECT 0.7350 0.8810 0.7850 1.0090 ;
        RECT 0.7350 0.8310 1.2410 0.8810 ;
        RECT 1.1910 0.8810 1.2410 1.5610 ;
    END
  END VSSG

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.1280 0.0300 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 2.1280 3.3740 ;
    END
  END VDD

  PIN VSS
    DIRECTION OUTPUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.1280 1.7020 ;
        RECT 1.3430 1.2010 1.3930 1.6420 ;
        RECT 1.0390 1.2010 1.0890 1.6420 ;
    END
  END VSS

  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0990 0.6700 1.3330 0.7300 ;
        RECT 1.1200 0.5530 1.3100 0.6700 ;
    END
    ANTENNAGATEAREA 0.0252 ;
  END SLEEP
  OBS
    LAYER NWELL ;
      RECT -0.1290 2.3510 2.2470 3.4520 ;
      RECT 0.2300 1.9040 1.8970 2.3510 ;
      RECT 0.2300 0.9930 0.4930 1.9040 ;
      RECT 1.6000 0.9930 1.8970 1.9040 ;
      RECT -0.1190 0.9160 0.4930 0.9930 ;
      RECT 1.6000 0.9160 2.2620 0.9930 ;
      RECT -0.1190 -0.1010 2.2620 0.9160 ;
    LAYER PO ;
      RECT 1.2770 2.0870 1.3070 3.1920 ;
      RECT 1.1250 2.0870 1.1550 3.1920 ;
      RECT 1.4290 2.0870 1.4590 3.1920 ;
      RECT 0.9730 2.0870 1.0030 3.1920 ;
      RECT 1.5810 2.0870 1.6110 3.1920 ;
      RECT 0.8210 2.0870 0.8510 3.1920 ;
      RECT 0.6690 2.0870 0.6990 3.1920 ;
      RECT 1.7330 2.0870 1.7630 3.1920 ;
      RECT 1.8850 2.0870 1.9150 3.1920 ;
      RECT 2.0370 2.0870 2.0670 3.1920 ;
      RECT 0.5170 2.0870 0.5470 3.1920 ;
      RECT 0.3650 2.0870 0.3950 3.1920 ;
      RECT 0.0610 2.0870 0.0910 3.1920 ;
      RECT 0.2130 2.0870 0.2430 3.1920 ;
      RECT 0.2130 0.5160 0.2430 1.6210 ;
      RECT 0.0610 0.5160 0.0910 1.6210 ;
      RECT 0.3650 0.5160 0.3950 1.6210 ;
      RECT 0.5170 0.5160 0.5470 1.6210 ;
      RECT 2.0370 0.5160 2.0670 1.6210 ;
      RECT 1.8850 0.5160 1.9150 1.6210 ;
      RECT 1.5810 0.5160 1.6110 1.6210 ;
      RECT 1.7330 0.5160 1.7630 1.6210 ;
      RECT 0.6690 0.5160 0.6990 1.6210 ;
      RECT 0.8210 0.5160 0.8510 1.6210 ;
      RECT 0.9730 0.5160 1.0030 1.6210 ;
      RECT 1.4290 0.5160 1.4590 1.6210 ;
      RECT 1.1250 0.5160 1.1550 1.6210 ;
      RECT 1.2770 0.5160 1.3070 1.6210 ;
  END
END FOOTX2_LVT

MACRO FOOTX32_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.688 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VSSG
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.6660 1.0090 0.8560 1.1190 ;
        RECT 0.7350 1.1190 0.7850 1.1650 ;
        RECT 0.7350 0.8810 0.7850 1.0090 ;
        RECT 0.7350 0.8310 5.8010 0.8810 ;
        RECT 3.3190 0.8810 3.3690 1.5610 ;
        RECT 3.6230 0.8810 3.6730 1.5610 ;
        RECT 3.9270 0.8810 3.9770 1.5610 ;
        RECT 4.2310 0.8810 4.2810 1.5610 ;
        RECT 4.5350 0.8810 4.5850 1.5610 ;
        RECT 4.8390 0.8810 4.8890 1.5610 ;
        RECT 5.1430 0.8810 5.1930 1.5610 ;
        RECT 5.4470 0.8810 5.4970 1.5610 ;
        RECT 2.1030 0.8810 2.1530 1.5610 ;
        RECT 2.4070 0.8810 2.4570 1.5610 ;
        RECT 2.7110 0.8810 2.7610 1.5610 ;
        RECT 3.0150 0.8810 3.0650 1.5610 ;
        RECT 1.7990 0.8810 1.8490 1.5610 ;
        RECT 1.4950 0.8810 1.5450 1.5610 ;
        RECT 5.7510 0.8810 5.8010 1.5610 ;
        RECT 1.1910 0.8810 1.2410 1.5610 ;
    END
  END VSSG

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 6.6880 0.0300 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 6.6880 3.3740 ;
    END
  END VDD

  PIN VSS
    DIRECTION OUTPUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 6.6880 1.7020 ;
        RECT 5.9030 1.2000 5.9530 1.6420 ;
        RECT 5.5990 1.2000 5.6490 1.6420 ;
        RECT 5.2950 1.2000 5.3450 1.6420 ;
        RECT 4.9910 1.2000 5.0410 1.6420 ;
        RECT 4.6870 1.2000 4.7370 1.6420 ;
        RECT 4.3830 1.2010 4.4330 1.6420 ;
        RECT 4.0790 1.2010 4.1290 1.6420 ;
        RECT 3.7750 1.2010 3.8250 1.6420 ;
        RECT 3.4710 1.2010 3.5210 1.6420 ;
        RECT 3.1670 1.2010 3.2170 1.6420 ;
        RECT 2.8630 1.2010 2.9130 1.6420 ;
        RECT 2.5590 1.2010 2.6090 1.6420 ;
        RECT 2.2550 1.2010 2.3050 1.6420 ;
        RECT 1.9510 1.2010 2.0010 1.6420 ;
        RECT 1.0390 1.2010 1.0890 1.6420 ;
        RECT 1.6470 1.2010 1.6970 1.6420 ;
        RECT 1.3430 1.2010 1.3930 1.6420 ;
    END
  END VSS

  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0990 0.6700 5.8930 0.7300 ;
        RECT 1.1200 0.5530 1.3100 0.6700 ;
    END
    ANTENNAGATEAREA 0.4032 ;
  END SLEEP
  OBS
    LAYER NWELL ;
      RECT -0.2050 2.3510 6.8540 3.5630 ;
      RECT 0.2300 1.6990 6.4580 2.3510 ;
      RECT 0.2300 0.9930 0.4910 1.6990 ;
      RECT 6.1750 0.9930 6.4580 1.6990 ;
      RECT -0.1390 0.6330 0.4910 0.9930 ;
      RECT 6.1750 0.6330 6.8520 0.9930 ;
      RECT -0.1390 -0.1700 6.8520 0.6330 ;
    LAYER PO ;
      RECT 5.2290 0.4870 5.2590 1.6210 ;
      RECT 5.3810 0.4870 5.4110 1.6210 ;
      RECT 5.5330 0.4870 5.5630 1.6210 ;
      RECT 5.6850 0.4870 5.7150 1.6210 ;
      RECT 5.9890 0.4870 6.0190 1.6210 ;
      RECT 5.8370 0.4870 5.8670 1.6210 ;
      RECT 2.4930 0.4870 2.5230 1.6210 ;
      RECT 2.6450 0.4870 2.6750 1.6210 ;
      RECT 2.7970 0.4870 2.8270 1.6210 ;
      RECT 2.9490 0.4870 2.9790 1.6210 ;
      RECT 3.1010 0.4870 3.1310 1.6210 ;
      RECT 3.2530 0.4870 3.2830 1.6210 ;
      RECT 3.4050 0.4870 3.4350 1.6210 ;
      RECT 3.5570 0.4870 3.5870 1.6210 ;
      RECT 2.0370 0.4870 2.0670 1.6210 ;
      RECT 0.6690 0.4870 0.6990 1.6210 ;
      RECT 2.1890 2.0380 2.2190 3.1720 ;
      RECT 1.5810 0.4870 1.6110 1.6210 ;
      RECT 0.8210 0.4870 0.8510 1.6210 ;
      RECT 6.1410 0.4870 6.1710 1.6210 ;
      RECT 0.9730 0.4870 1.0030 1.6210 ;
      RECT 1.4290 0.4870 1.4590 1.6210 ;
      RECT 1.7330 0.4870 1.7630 1.6210 ;
      RECT 1.1250 0.4870 1.1550 1.6210 ;
      RECT 2.3410 0.4870 2.3710 1.6210 ;
      RECT 1.8850 2.0380 1.9150 3.1720 ;
      RECT 1.2770 0.4870 1.3070 1.6210 ;
      RECT 2.1890 0.4870 2.2190 1.6210 ;
      RECT 1.8850 0.4870 1.9150 1.6210 ;
      RECT 6.4450 0.4870 6.4750 1.6210 ;
      RECT 6.5970 0.4870 6.6270 1.6210 ;
      RECT 6.2930 0.4870 6.3230 1.6210 ;
      RECT 0.0610 0.4870 0.0910 1.6210 ;
      RECT 0.5170 0.4870 0.5470 1.6210 ;
      RECT 0.3650 0.4870 0.3950 1.6210 ;
      RECT 0.2130 0.4870 0.2430 1.6210 ;
      RECT 6.4450 2.0380 6.4750 3.1720 ;
      RECT 6.5970 2.0380 6.6270 3.1720 ;
      RECT 6.2930 2.0380 6.3230 3.1720 ;
      RECT 0.0610 2.0380 0.0910 3.1720 ;
      RECT 0.5170 2.0380 0.5470 3.1720 ;
      RECT 0.3650 2.0380 0.3950 3.1720 ;
      RECT 0.2130 2.0380 0.2430 3.1720 ;
      RECT 3.7090 2.0380 3.7390 3.1720 ;
      RECT 3.8610 2.0380 3.8910 3.1720 ;
      RECT 4.0130 2.0380 4.0430 3.1720 ;
      RECT 4.1650 2.0380 4.1950 3.1720 ;
      RECT 4.3170 2.0380 4.3470 3.1720 ;
      RECT 4.4690 2.0380 4.4990 3.1720 ;
      RECT 4.6210 2.0380 4.6510 3.1720 ;
      RECT 4.7730 2.0380 4.8030 3.1720 ;
      RECT 4.9250 2.0380 4.9550 3.1720 ;
      RECT 5.0770 2.0380 5.1070 3.1720 ;
      RECT 5.2290 2.0380 5.2590 3.1720 ;
      RECT 5.3810 2.0380 5.4110 3.1720 ;
      RECT 5.5330 2.0380 5.5630 3.1720 ;
      RECT 5.6850 2.0380 5.7150 3.1720 ;
      RECT 5.9890 2.0380 6.0190 3.1720 ;
      RECT 5.8370 2.0380 5.8670 3.1720 ;
      RECT 2.4930 2.0380 2.5230 3.1720 ;
      RECT 2.6450 2.0380 2.6750 3.1720 ;
      RECT 2.7970 2.0380 2.8270 3.1720 ;
      RECT 2.9490 2.0380 2.9790 3.1720 ;
      RECT 3.1010 2.0380 3.1310 3.1720 ;
      RECT 3.2530 2.0380 3.2830 3.1720 ;
      RECT 3.4050 2.0380 3.4350 3.1720 ;
      RECT 3.5570 2.0380 3.5870 3.1720 ;
      RECT 2.0370 2.0380 2.0670 3.1720 ;
      RECT 0.6690 2.0380 0.6990 3.1720 ;
      RECT 1.5810 2.0380 1.6110 3.1720 ;
      RECT 0.8210 2.0380 0.8510 3.1720 ;
      RECT 6.1410 2.0380 6.1710 3.1720 ;
      RECT 0.9730 2.0380 1.0030 3.1720 ;
      RECT 1.4290 2.0380 1.4590 3.1720 ;
      RECT 1.7330 2.0380 1.7630 3.1720 ;
      RECT 1.1250 2.0380 1.1550 3.1720 ;
      RECT 2.3410 2.0380 2.3710 3.1720 ;
      RECT 1.2770 2.0380 1.3070 3.1720 ;
      RECT 3.7090 0.4870 3.7390 1.6210 ;
      RECT 3.8610 0.4870 3.8910 1.6210 ;
      RECT 4.0130 0.4870 4.0430 1.6210 ;
      RECT 4.1650 0.4870 4.1950 1.6210 ;
      RECT 4.3170 0.4870 4.3470 1.6210 ;
      RECT 4.4690 0.4870 4.4990 1.6210 ;
      RECT 4.6210 0.4870 4.6510 1.6210 ;
      RECT 4.7730 0.4870 4.8030 1.6210 ;
      RECT 4.9250 0.4870 4.9550 1.6210 ;
      RECT 5.0770 0.4870 5.1070 1.6210 ;
  END
END FOOTX32_LVT

MACRO FOOTX4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.28 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VSSG
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.5140 1.0090 0.7040 1.1190 ;
        RECT 0.5830 1.1190 0.6330 1.1650 ;
        RECT 0.5830 0.8810 0.6330 1.0090 ;
        RECT 0.5830 0.8310 1.3930 0.8810 ;
        RECT 1.3430 0.8810 1.3930 1.5610 ;
        RECT 1.0390 0.8810 1.0890 1.5610 ;
    END
  END VSSG

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.2800 0.0300 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 2.2800 3.3740 ;
    END
  END VDD

  PIN VSS
    DIRECTION OUTPUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.2800 1.7020 ;
        RECT 0.8870 1.2010 0.9370 1.6420 ;
        RECT 1.4950 1.2010 1.5450 1.6420 ;
        RECT 1.1910 1.2010 1.2410 1.6420 ;
    END
  END VSS

  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9470 0.6700 1.4850 0.7300 ;
        RECT 0.9680 0.5530 1.1580 0.6700 ;
    END
    ANTENNAGATEAREA 0.0504 ;
  END SLEEP
  OBS
    LAYER NWELL ;
      RECT -0.0820 2.3510 2.3550 3.4480 ;
      RECT 0.2310 1.6890 1.9520 2.3510 ;
      RECT 0.2310 0.9930 0.4660 1.6890 ;
      RECT 1.6400 0.9930 1.9520 1.6890 ;
      RECT -0.0800 0.8150 0.4660 0.9930 ;
      RECT 1.6400 0.8150 2.3840 0.9930 ;
      RECT -0.0800 -0.1150 2.3840 0.8150 ;
    LAYER PO ;
      RECT 1.1250 2.0450 1.1550 3.1790 ;
      RECT 0.9730 2.0450 1.0030 3.1790 ;
      RECT 1.5810 2.0450 1.6110 3.1790 ;
      RECT 1.2770 2.0450 1.3070 3.1790 ;
      RECT 0.8210 2.0450 0.8510 3.1790 ;
      RECT 1.7330 2.0450 1.7630 3.1790 ;
      RECT 0.6690 2.0450 0.6990 3.1790 ;
      RECT 0.0610 2.0450 0.0910 3.1790 ;
      RECT 2.0370 0.4870 2.0670 1.6210 ;
      RECT 1.7330 0.4870 1.7630 1.6210 ;
      RECT 0.2130 2.0450 0.2430 3.1790 ;
      RECT 1.8850 0.4870 1.9150 1.6210 ;
      RECT 0.0610 0.4870 0.0910 1.6210 ;
      RECT 0.2130 0.4870 0.2430 1.6210 ;
      RECT 0.5170 0.4870 0.5470 1.6210 ;
      RECT 0.6690 0.4870 0.6990 1.6210 ;
      RECT 2.1890 2.0450 2.2190 3.1790 ;
      RECT 0.3650 0.4870 0.3950 1.6210 ;
      RECT 2.1890 0.4870 2.2190 1.6210 ;
      RECT 0.5170 2.0450 0.5470 3.1790 ;
      RECT 2.0370 2.0450 2.0670 3.1790 ;
      RECT 0.3650 2.0450 0.3950 3.1790 ;
      RECT 1.8850 2.0450 1.9150 3.1790 ;
      RECT 1.4290 0.4870 1.4590 1.6210 ;
      RECT 0.8210 0.4870 0.8510 1.6210 ;
      RECT 1.2770 0.4870 1.3070 1.6210 ;
      RECT 1.5810 0.4870 1.6110 1.6210 ;
      RECT 0.9730 0.4870 1.0030 1.6210 ;
      RECT 1.1250 0.4870 1.1550 1.6210 ;
      RECT 1.4290 2.0450 1.4590 3.1790 ;
  END
END FOOTX4_LVT

MACRO FOOTX8_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.04 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VSSG
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.6660 1.0090 0.8560 1.1190 ;
        RECT 0.7350 1.1190 0.7850 1.1650 ;
        RECT 0.7350 0.8810 0.7850 1.0090 ;
        RECT 0.7350 0.8310 2.1530 0.8810 ;
        RECT 1.7990 0.8810 1.8490 1.5610 ;
        RECT 1.4950 0.8810 1.5450 1.5610 ;
        RECT 2.1030 0.8810 2.1530 1.5610 ;
        RECT 1.1910 0.8810 1.2410 1.5610 ;
    END
  END VSSG

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.0400 0.0300 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 3.0400 3.3740 ;
    END
  END VDD

  PIN VSS
    DIRECTION OUTPUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.0400 1.7020 ;
        RECT 2.2550 1.2010 2.3050 1.6420 ;
        RECT 1.9510 1.2010 2.0010 1.6420 ;
        RECT 1.0390 1.2010 1.0890 1.6420 ;
        RECT 1.6470 1.2010 1.6970 1.6420 ;
        RECT 1.3430 1.2010 1.3930 1.6420 ;
    END
  END VSS

  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0990 0.6700 2.2450 0.7300 ;
        RECT 1.1200 0.5530 1.3100 0.6700 ;
    END
    ANTENNAGATEAREA 0.1008 ;
  END SLEEP
  OBS
    LAYER NWELL ;
      RECT -0.1330 2.3510 3.1600 3.5180 ;
      RECT 0.2320 1.6540 2.8060 2.3510 ;
      RECT 0.2320 0.9930 0.5760 1.6540 ;
      RECT 2.4580 0.9930 2.8060 1.6540 ;
      RECT -0.1270 0.7800 0.5760 0.9930 ;
      RECT 2.4580 0.7800 3.1460 0.9930 ;
      RECT -0.1270 -0.1750 3.1460 0.7800 ;
    LAYER PO ;
      RECT 1.8850 2.0590 1.9150 3.1930 ;
      RECT 2.1890 2.0590 2.2190 3.1930 ;
      RECT 1.2770 2.0590 1.3070 3.1930 ;
      RECT 2.3410 2.0590 2.3710 3.1930 ;
      RECT 1.1250 2.0590 1.1550 3.1930 ;
      RECT 1.7330 2.0590 1.7630 3.1930 ;
      RECT 1.4290 2.0590 1.4590 3.1930 ;
      RECT 0.9730 2.0590 1.0030 3.1930 ;
      RECT 2.4930 2.0590 2.5230 3.1930 ;
      RECT 0.8210 2.0590 0.8510 3.1930 ;
      RECT 1.5810 2.0590 1.6110 3.1930 ;
      RECT 0.6690 2.0590 0.6990 3.1930 ;
      RECT 2.0370 2.0590 2.0670 3.1930 ;
      RECT 2.7970 2.0590 2.8270 3.1930 ;
      RECT 2.9490 2.0590 2.9790 3.1930 ;
      RECT 2.6450 2.0590 2.6750 3.1930 ;
      RECT 0.0610 2.0590 0.0910 3.1930 ;
      RECT 0.2130 2.0590 0.2430 3.1930 ;
      RECT 0.5170 2.0590 0.5470 3.1930 ;
      RECT 0.3650 2.0590 0.3950 3.1930 ;
      RECT 0.2130 0.1520 0.2430 1.6210 ;
      RECT 0.3650 0.1520 0.3950 1.6210 ;
      RECT 0.6690 0.1520 0.6990 1.6210 ;
      RECT 0.5170 0.1520 0.5470 1.6210 ;
      RECT 0.0610 0.1520 0.0910 1.6210 ;
      RECT 2.7970 0.1520 2.8270 1.6210 ;
      RECT 2.9490 0.1520 2.9790 1.6210 ;
      RECT 2.6450 0.1520 2.6750 1.6210 ;
      RECT 2.0370 0.1520 2.0670 1.6210 ;
      RECT 1.5810 0.1520 1.6110 1.6210 ;
      RECT 0.8210 0.1520 0.8510 1.6210 ;
      RECT 2.4930 0.1520 2.5230 1.6210 ;
      RECT 0.9730 0.1520 1.0030 1.6210 ;
      RECT 1.4290 0.1520 1.4590 1.6210 ;
      RECT 1.7330 0.1520 1.7630 1.6210 ;
      RECT 1.1250 0.1520 1.1550 1.6210 ;
      RECT 2.3410 0.1520 2.3710 1.6210 ;
      RECT 1.2770 0.1520 1.3070 1.6210 ;
      RECT 2.1890 0.1520 2.2190 1.6210 ;
      RECT 1.8850 0.1520 1.9150 1.6210 ;
  END
END FOOTX8_LVT

MACRO HADDX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.976 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6310 0.1380 1.7210 0.1880 ;
        RECT 1.6710 0.1880 1.7210 0.8480 ;
        RECT 1.6710 0.8480 1.8790 0.9100 ;
        RECT 1.6310 0.9100 1.8790 0.9580 ;
        RECT 1.6310 0.9580 1.7210 0.9600 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END SO

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5070 0.6030 1.1650 0.6530 ;
        RECT 0.5070 0.5520 0.5570 0.6030 ;
        RECT 0.6490 0.6530 0.8150 0.6630 ;
        RECT 0.6490 0.5530 0.8150 0.6030 ;
        RECT 1.1150 0.5150 1.1650 0.6030 ;
    END
    ANTENNAGATEAREA 0.0513 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.7460 1.0290 0.7960 ;
        RECT 0.3450 0.7960 0.5110 0.8150 ;
        RECT 0.3450 0.7050 0.5110 0.7460 ;
    END
    ANTENNAGATEAREA 0.0513 ;
  END A0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.9760 1.7020 ;
        RECT 1.0390 1.3180 1.0890 1.6420 ;
        RECT 1.4950 1.3420 1.5450 1.6420 ;
        RECT 0.2790 1.3230 0.3290 1.6420 ;
        RECT 0.7350 1.3230 0.7850 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.9760 0.0300 ;
        RECT 0.7350 0.0300 0.7850 0.2540 ;
        RECT 0.8870 0.0300 0.9370 0.2610 ;
        RECT 1.4950 0.0300 1.5450 0.1370 ;
        RECT 1.4790 0.1370 1.5610 0.1870 ;
    END
  END VSS

  PIN C1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3150 0.5610 1.3650 1.0000 ;
        RECT 1.3150 1.0000 1.5750 1.1190 ;
        RECT 1.3150 0.4740 1.3930 0.5610 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END C1
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 2.0910 1.7730 ;
    LAYER M1 ;
      RECT 1.4520 0.3870 1.5020 0.6130 ;
      RECT 1.4190 0.6130 1.5020 0.6630 ;
      RECT 1.1750 0.3370 1.5020 0.3870 ;
      RECT 1.4190 0.6630 1.4690 0.7360 ;
      RECT 1.2150 1.1760 1.2650 1.3170 ;
      RECT 1.1910 1.3170 1.2650 1.4110 ;
      RECT 0.8110 1.1260 1.2650 1.1760 ;
      RECT 1.2150 0.3870 1.2650 1.1260 ;
      RECT 0.8110 0.9390 0.8610 1.1260 ;
      RECT 0.6380 0.8890 0.8610 0.9390 ;
      RECT 0.2630 0.1740 0.6550 0.2240 ;
      RECT 1.5710 0.2870 1.6210 0.7340 ;
      RECT 1.0130 0.2380 1.6210 0.2870 ;
      RECT 1.0130 0.2370 1.5810 0.2380 ;
      RECT 1.0130 0.2870 1.0630 0.3600 ;
      RECT 0.2390 0.3600 1.0630 0.4100 ;
      RECT 0.2390 1.0570 0.6490 1.1070 ;
      RECT 0.2390 0.4100 0.2890 1.0570 ;
    LAYER PO ;
      RECT 0.3650 0.0710 0.3950 1.6090 ;
      RECT 0.5170 0.0710 0.5470 1.6090 ;
      RECT 0.9730 0.0710 1.0030 1.6090 ;
      RECT 1.5810 0.0710 1.6110 1.6160 ;
      RECT 1.2770 0.0710 1.3070 1.6090 ;
      RECT 0.0610 0.0710 0.0910 1.6090 ;
      RECT 1.1250 0.0710 1.1550 1.6090 ;
      RECT 0.8210 0.0670 0.8510 1.6090 ;
      RECT 1.4290 0.0710 1.4590 1.6160 ;
      RECT 0.2130 0.0710 0.2430 1.6090 ;
      RECT 0.6690 0.0710 0.6990 1.6090 ;
      RECT 1.8850 0.0710 1.9150 1.6090 ;
      RECT 1.7330 0.0710 1.7630 1.6090 ;
  END
END HADDX1_LVT

MACRO HADDX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.28 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7980 0.3050 1.8480 0.3250 ;
        RECT 1.7980 0.3250 2.0670 0.3750 ;
        RECT 2.0170 0.3750 2.0670 0.9570 ;
        RECT 1.7980 0.3750 1.8480 0.3960 ;
        RECT 2.0170 0.9570 2.1830 1.0170 ;
        RECT 1.7830 1.0170 2.1830 1.0670 ;
        RECT 2.0170 1.0670 2.1830 1.1190 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END SO

  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4850 0.5870 1.1640 0.6370 ;
        RECT 0.5530 0.6370 0.6630 0.6630 ;
        RECT 0.5530 0.5530 0.6630 0.5870 ;
        RECT 1.1140 0.6370 1.1640 0.6530 ;
        RECT 1.1140 0.5710 1.1640 0.5870 ;
    END
    ANTENNAGATEAREA 0.0513 ;
  END B0

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3390 0.7130 1.0290 0.7630 ;
        RECT 0.3450 0.7630 0.5110 0.8150 ;
        RECT 0.3450 0.7050 0.5110 0.7130 ;
    END
    ANTENNAGATEAREA 0.0513 ;
  END A0

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.2800 1.7020 ;
        RECT 1.0390 1.3190 1.0890 1.6420 ;
        RECT 1.3430 1.3630 1.3930 1.6420 ;
        RECT 1.6470 1.3630 1.6970 1.6420 ;
        RECT 1.9510 1.3630 2.0010 1.6420 ;
        RECT 0.2790 1.3190 0.3290 1.6420 ;
        RECT 0.7350 1.3190 0.7850 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.2800 0.0300 ;
        RECT 0.7350 0.0300 0.7850 0.2540 ;
        RECT 0.8870 0.0300 0.9370 0.2590 ;
        RECT 1.9510 0.0300 2.0010 0.2100 ;
        RECT 1.3430 0.0300 1.3930 0.1370 ;
        RECT 1.6470 0.0300 1.6970 0.1370 ;
        RECT 1.3270 0.1370 1.4090 0.1870 ;
        RECT 1.6310 0.1370 1.7130 0.1870 ;
    END
  END VSS

  PIN C1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3150 0.5450 1.3650 1.1610 ;
        RECT 1.3150 1.1610 1.5750 1.2940 ;
        RECT 1.3150 0.4950 1.5450 0.5450 ;
        RECT 1.4950 0.5450 1.5450 0.5610 ;
        RECT 1.4950 0.4740 1.5450 0.4950 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END C1
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 2.3950 1.7730 ;
    LAYER M1 ;
      RECT 1.1750 0.3370 1.6450 0.3870 ;
      RECT 1.4190 0.6390 1.6450 0.7270 ;
      RECT 1.5950 0.7270 1.6450 0.7290 ;
      RECT 1.5950 0.3870 1.6450 0.6390 ;
      RECT 0.8110 0.9390 0.8610 1.1260 ;
      RECT 0.6380 0.8890 0.8610 0.9390 ;
      RECT 0.8110 1.1260 1.2650 1.1760 ;
      RECT 1.2150 1.1760 1.2650 1.3170 ;
      RECT 1.1910 1.3170 1.2650 1.4110 ;
      RECT 1.2150 0.3870 1.2650 1.1260 ;
      RECT 1.6950 0.6390 1.9290 0.7270 ;
      RECT 1.6950 0.7270 1.7450 0.7300 ;
      RECT 1.6950 0.2870 1.7450 0.6390 ;
      RECT 1.0130 0.2370 1.7450 0.2870 ;
      RECT 0.2390 1.0570 0.6490 1.1070 ;
      RECT 0.2390 0.3590 0.2890 1.0570 ;
      RECT 1.0130 0.2870 1.0630 0.3090 ;
      RECT 0.2390 0.3090 1.0630 0.3590 ;
      RECT 0.2630 0.1700 0.6550 0.2200 ;
    LAYER PO ;
      RECT 2.0370 0.0710 2.0670 1.6090 ;
      RECT 2.1890 0.0710 2.2190 1.6090 ;
      RECT 0.3650 0.0710 0.3950 1.6090 ;
      RECT 0.5170 0.0710 0.5470 1.6090 ;
      RECT 0.9730 0.0710 1.0030 1.6090 ;
      RECT 1.5810 0.0710 1.6110 1.6090 ;
      RECT 1.2770 0.0710 1.3070 1.6090 ;
      RECT 0.0610 0.0710 0.0910 1.6090 ;
      RECT 1.1250 0.0710 1.1550 1.6090 ;
      RECT 0.8210 0.0670 0.8510 1.6090 ;
      RECT 1.4290 0.0710 1.4590 1.6090 ;
      RECT 0.2130 0.0710 0.2430 1.6090 ;
      RECT 0.6690 0.0710 0.6990 1.6090 ;
      RECT 1.8850 0.0710 1.9150 1.6090 ;
      RECT 1.7330 0.0710 1.7630 1.6090 ;
  END
END HADDX2_LVT

MACRO HEAD2X16_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.56 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SLEEPOUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6470 0.8060 3.8150 0.8660 ;
        RECT 1.6470 0.7950 1.6970 0.8060 ;
        RECT 3.4710 0.8660 3.5210 1.3580 ;
        RECT 3.4710 0.7950 3.5210 0.8060 ;
        RECT 3.1670 0.8660 3.2170 1.3580 ;
        RECT 3.1670 0.7950 3.2170 0.8060 ;
        RECT 2.8630 0.8660 2.9130 1.3580 ;
        RECT 2.8630 0.7950 2.9130 0.8060 ;
        RECT 2.5590 0.8660 2.6090 1.3580 ;
        RECT 2.5590 0.7950 2.6090 0.8060 ;
        RECT 2.2550 0.8660 2.3050 1.3580 ;
        RECT 2.2550 0.7950 2.3050 0.8060 ;
        RECT 1.9510 0.8660 2.0010 1.3580 ;
        RECT 1.9510 0.7950 2.0010 0.8060 ;
        RECT 3.7650 0.6630 3.8150 0.8060 ;
        RECT 1.6470 0.8660 1.6970 1.0840 ;
        RECT 3.7320 0.5620 3.8550 0.6630 ;
        RECT 1.3270 1.0840 1.6970 1.1440 ;
        RECT 1.3430 0.5520 3.8550 0.5620 ;
        RECT 1.3430 1.1440 1.3930 1.3580 ;
        RECT 1.3430 1.0730 1.3930 1.0840 ;
        RECT 1.6470 1.1440 1.6970 1.3580 ;
        RECT 1.3430 0.5020 3.8510 0.5520 ;
        RECT 1.3430 0.1800 1.3930 0.5020 ;
        RECT 3.4710 0.1790 3.5210 0.5020 ;
        RECT 3.1670 0.1790 3.2170 0.5020 ;
        RECT 2.8630 0.1790 2.9130 0.5020 ;
        RECT 2.5590 0.1790 2.6090 0.5020 ;
        RECT 2.2550 0.1790 2.3050 0.5020 ;
        RECT 1.9510 0.1800 2.0010 0.5020 ;
        RECT 1.6470 0.1800 1.6970 0.5020 ;
    END
    ANTENNADIFFAREA 1.1904 ;
  END SLEEPOUT

  PIN VDDG
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 3.5520 2.0730 3.7420 2.1830 ;
        RECT 3.6180 2.0110 3.6780 2.0730 ;
        RECT 3.6180 2.1830 3.6780 2.4930 ;
        RECT 1.0380 2.4930 3.9170 2.5430 ;
        RECT 1.9510 1.8370 2.0010 2.4930 ;
        RECT 1.6470 1.8370 1.6970 2.4930 ;
        RECT 1.3430 1.8370 1.3930 2.4930 ;
        RECT 1.0390 1.8370 1.0890 2.4930 ;
        RECT 3.1670 1.8370 3.2170 2.4930 ;
        RECT 2.8630 1.8370 2.9130 2.4930 ;
        RECT 2.5590 1.8370 2.6090 2.4930 ;
        RECT 2.2550 1.8370 2.3050 2.4930 ;
    END
  END VDDG

  PIN VDD
    DIRECTION OUTPUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.5600 1.7020 ;
        RECT 3.3190 1.7020 3.3690 2.3090 ;
        RECT 3.0150 1.7020 3.0650 2.3090 ;
        RECT 2.7110 1.7020 2.7610 2.3090 ;
        RECT 2.4070 1.7020 2.4570 2.3100 ;
        RECT 2.1030 1.7020 2.1530 2.3100 ;
        RECT 1.7990 1.7020 1.8490 2.3100 ;
        RECT 1.4950 1.7020 1.5450 2.3100 ;
        RECT 0.8870 1.7020 0.9370 2.4940 ;
        RECT 1.1910 1.7020 1.2410 2.3100 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.5600 0.0300 ;
        RECT 3.6230 0.0300 3.6730 0.3820 ;
        RECT 3.3190 0.0300 3.3690 0.3820 ;
        RECT 3.0150 0.0300 3.0650 0.3820 ;
        RECT 2.7110 0.0300 2.7610 0.3820 ;
        RECT 2.4070 0.0300 2.4570 0.3820 ;
        RECT 2.1030 0.0300 2.1530 0.3820 ;
        RECT 1.7990 0.0300 1.8490 0.3820 ;
        RECT 1.1910 0.0300 1.2410 0.5660 ;
        RECT 1.4950 0.0300 1.5450 0.3820 ;
        RECT 0.8870 0.0300 0.9370 0.3820 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 4.5600 3.3740 ;
    END
  END VSS

  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7950 0.6570 1.1810 0.7170 ;
        RECT 0.8310 0.7170 0.9910 0.8150 ;
    END
    ANTENNAGATEAREA 0.1098 ;
  END SLEEP
  OBS
    LAYER NWELL ;
      RECT 0.5710 0.6790 3.9810 2.6650 ;
    LAYER M1 ;
      RECT 0.8870 1.4590 3.9170 1.5190 ;
      RECT 3.6230 1.0480 3.6730 1.4590 ;
      RECT 1.1910 1.0480 1.2410 1.4590 ;
      RECT 0.8870 1.0480 0.9370 1.4590 ;
      RECT 1.4950 1.2340 1.5450 1.4590 ;
      RECT 1.7990 1.0480 1.8490 1.4590 ;
      RECT 2.1030 1.0480 2.1530 1.4590 ;
      RECT 2.4070 1.0480 2.4570 1.4590 ;
      RECT 2.7110 1.0480 2.7610 1.4590 ;
      RECT 3.0150 1.0480 3.0650 1.4590 ;
      RECT 3.3190 1.0480 3.3690 1.4590 ;
      RECT 1.2510 0.6560 3.6130 0.7160 ;
      RECT 0.7350 0.9900 0.7850 1.3580 ;
      RECT 0.7350 0.1800 0.7850 0.5020 ;
      RECT 1.0390 0.9900 1.0890 1.3580 ;
      RECT 0.6590 0.5020 1.0890 0.5620 ;
      RECT 1.0390 0.1800 1.0890 0.5020 ;
      RECT 1.2510 0.7160 1.3010 0.9300 ;
      RECT 0.6590 0.9300 1.3010 0.9900 ;
      RECT 0.6590 0.5620 0.7090 0.9300 ;
      RECT 0.6430 2.6030 3.3090 2.6530 ;
    LAYER PO ;
      RECT 1.7330 0.1200 1.7630 1.6070 ;
      RECT 2.0370 1.7070 2.0670 3.2630 ;
      RECT 2.1890 1.7070 2.2190 3.2630 ;
      RECT 3.8610 0.1200 3.8910 3.2630 ;
      RECT 2.0370 0.1200 2.0670 1.6070 ;
      RECT 1.7330 1.7070 1.7630 3.2630 ;
      RECT 0.6690 0.1200 0.6990 3.2630 ;
      RECT 0.9730 1.7070 1.0030 3.2630 ;
      RECT 1.5810 1.7070 1.6110 3.2630 ;
      RECT 1.4290 1.7070 1.4590 3.2630 ;
      RECT 0.8210 1.7070 0.8510 3.2630 ;
      RECT 0.8210 0.1190 0.8510 1.6070 ;
      RECT 1.1250 1.7070 1.1550 3.2630 ;
      RECT 1.5810 0.1200 1.6110 1.6070 ;
      RECT 3.5570 1.7070 3.5870 3.2630 ;
      RECT 0.9730 0.1200 1.0030 1.6070 ;
      RECT 1.4290 0.1200 1.4590 1.6070 ;
      RECT 1.1250 0.1200 1.1550 1.6070 ;
      RECT 1.2770 0.1200 1.3070 1.6070 ;
      RECT 1.2770 1.7070 1.3070 3.2630 ;
      RECT 4.4690 1.7070 4.4990 3.2630 ;
      RECT 4.3170 1.7070 4.3470 3.2630 ;
      RECT 4.0130 1.7070 4.0430 3.2590 ;
      RECT 4.1650 1.7070 4.1950 3.2590 ;
      RECT 4.1650 0.1200 4.1950 1.6070 ;
      RECT 4.3170 0.1200 4.3470 1.6070 ;
      RECT 4.4690 0.1200 4.4990 1.6070 ;
      RECT 4.0130 0.1200 4.0430 1.6070 ;
      RECT 0.0610 0.1190 0.0910 1.6070 ;
      RECT 0.2130 0.1200 0.2430 1.6070 ;
      RECT 0.3650 0.1200 0.3950 1.6070 ;
      RECT 0.5170 0.1200 0.5470 1.6070 ;
      RECT 0.2130 1.7070 0.2430 3.2630 ;
      RECT 0.0610 1.7070 0.0910 3.2630 ;
      RECT 0.3650 1.7070 0.3950 3.2630 ;
      RECT 0.5170 1.7070 0.5470 3.2630 ;
      RECT 2.3410 1.7070 2.3710 3.2590 ;
      RECT 2.4930 1.7070 2.5230 3.2590 ;
      RECT 2.6450 1.7070 2.6750 3.2590 ;
      RECT 2.7970 1.7070 2.8270 3.2590 ;
      RECT 2.9490 1.7070 2.9790 3.2590 ;
      RECT 3.1010 1.7070 3.1310 3.2590 ;
      RECT 3.2530 1.7070 3.2830 3.2590 ;
      RECT 3.4050 1.7070 3.4350 3.2590 ;
      RECT 3.1010 0.1200 3.1310 1.6070 ;
      RECT 2.9490 0.1200 2.9790 1.6070 ;
      RECT 2.7970 0.1200 2.8270 1.6070 ;
      RECT 2.6450 0.1200 2.6750 1.6070 ;
      RECT 3.2530 0.1200 3.2830 1.6070 ;
      RECT 3.4050 0.1200 3.4350 1.6070 ;
      RECT 3.5570 0.1200 3.5870 1.6070 ;
      RECT 3.7090 0.1200 3.7390 1.6070 ;
      RECT 3.7090 1.7070 3.7390 3.2630 ;
      RECT 2.4930 0.1200 2.5230 1.6070 ;
      RECT 2.1890 0.1200 2.2190 1.6070 ;
      RECT 1.8850 1.7070 1.9150 3.2630 ;
      RECT 1.8850 0.1200 1.9150 1.6070 ;
      RECT 2.3410 0.1200 2.3710 1.6070 ;
  END
END HEAD2X16_LVT

MACRO HEAD2X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.28 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SLEEPOUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1910 1.0830 1.5210 1.1430 ;
        RECT 1.1910 1.1430 1.2410 1.4090 ;
        RECT 1.4710 0.6630 1.5210 1.0830 ;
        RECT 1.4520 0.5620 1.5750 0.6630 ;
        RECT 1.1910 0.5520 1.5750 0.5620 ;
        RECT 1.1910 0.5020 1.5710 0.5520 ;
        RECT 1.1910 0.1800 1.2410 0.5020 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END SLEEPOUT

  PIN VDDG
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 1.2720 2.0730 1.4620 2.1830 ;
        RECT 1.3380 2.0270 1.3980 2.0730 ;
        RECT 1.3380 2.1830 1.3980 2.4930 ;
        RECT 0.8860 2.4930 1.6370 2.5430 ;
        RECT 1.3380 2.5430 1.3980 2.5590 ;
        RECT 0.8870 1.8370 0.9370 2.4930 ;
    END
  END VDDG

  PIN VDD
    DIRECTION OUTPUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0300 1.6420 2.3100 1.7020 ;
        RECT 0.7350 1.7020 0.7850 2.4960 ;
        RECT 1.0390 1.7020 1.0890 2.4040 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.2800 0.0300 ;
        RECT 1.0390 0.0300 1.0890 0.5660 ;
        RECT 1.3430 0.0300 1.3930 0.3820 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 2.2800 3.3740 ;
    END
  END VSS

  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8530 0.7050 1.0130 0.8150 ;
        RECT 0.9630 0.6450 1.0130 0.7050 ;
    END
    ANTENNAGATEAREA 0.0366 ;
  END SLEEP
  OBS
    LAYER NWELL ;
      RECT 0.5710 0.6790 1.6730 2.6650 ;
      RECT 1.0800 1.9230 1.0830 1.9340 ;
    LAYER M1 ;
      RECT 1.0990 0.6560 1.3330 0.7160 ;
      RECT 0.8870 1.0160 0.9370 1.5190 ;
      RECT 0.6590 0.5020 0.9370 0.5620 ;
      RECT 0.8870 0.1800 0.9370 0.5020 ;
      RECT 1.1150 0.7160 1.1650 0.9560 ;
      RECT 0.6590 0.9560 1.1650 1.0160 ;
      RECT 0.6590 0.5620 0.7090 0.9560 ;
      RECT 1.3430 1.2340 1.3930 1.4590 ;
      RECT 1.0390 1.4590 1.6370 1.5190 ;
      RECT 1.0390 1.2340 1.0890 1.4590 ;
      RECT 0.6430 2.6030 1.0290 2.6530 ;
    LAYER PO ;
      RECT 2.1890 1.7070 2.2190 3.2180 ;
      RECT 1.7330 0.1150 1.7630 1.6070 ;
      RECT 1.8850 0.1150 1.9150 1.6070 ;
      RECT 2.0370 0.1150 2.0670 1.6070 ;
      RECT 0.0610 0.1150 0.0910 1.6070 ;
      RECT 0.2130 0.1150 0.2430 1.6070 ;
      RECT 0.3650 0.1150 0.3950 1.6070 ;
      RECT 1.7330 1.7070 1.7630 3.2180 ;
      RECT 1.8850 1.7070 1.9150 3.2180 ;
      RECT 0.0610 1.7070 0.0910 3.2180 ;
      RECT 2.0370 1.7070 2.0670 3.2180 ;
      RECT 0.2130 1.7070 0.2430 3.2180 ;
      RECT 1.5810 0.1200 1.6110 3.2150 ;
      RECT 0.5170 0.1200 0.5470 1.6070 ;
      RECT 0.8210 1.7070 0.8510 3.2180 ;
      RECT 1.4290 1.7210 1.4590 3.2150 ;
      RECT 1.2770 1.7210 1.3070 3.2150 ;
      RECT 0.3650 1.7070 0.3950 3.2180 ;
      RECT 0.6690 0.1190 0.6990 3.2180 ;
      RECT 0.9730 1.7070 1.0030 3.2180 ;
      RECT 1.4290 0.1200 1.4590 1.6210 ;
      RECT 0.8210 0.1200 0.8510 1.6070 ;
      RECT 1.2770 0.1200 1.3070 1.6210 ;
      RECT 0.5170 1.7070 0.5470 3.2090 ;
      RECT 0.9730 0.1200 1.0030 1.6070 ;
      RECT 1.1250 0.1200 1.1550 1.6210 ;
      RECT 1.1250 1.7210 1.1550 3.2180 ;
  END
END HEAD2X2_LVT

MACRO HEAD2X32_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.296 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 7.2960 0.0300 ;
        RECT 6.3590 0.0300 6.4090 0.3820 ;
        RECT 6.0550 0.0300 6.1050 0.3820 ;
        RECT 5.7510 0.0300 5.8010 0.3820 ;
        RECT 5.4470 0.0300 5.4970 0.3820 ;
        RECT 5.1430 0.0300 5.1930 0.3820 ;
        RECT 4.8390 0.0300 4.8890 0.3820 ;
        RECT 4.5350 0.0300 4.5850 0.3820 ;
        RECT 4.2310 0.0300 4.2810 0.3820 ;
        RECT 3.9270 0.0300 3.9770 0.3820 ;
        RECT 3.6230 0.0300 3.6730 0.3820 ;
        RECT 3.3190 0.0300 3.3690 0.3820 ;
        RECT 3.0150 0.0300 3.0650 0.3820 ;
        RECT 2.7110 0.0300 2.7610 0.3820 ;
        RECT 2.4070 0.0300 2.4570 0.3820 ;
        RECT 2.1030 0.0300 2.1530 0.3820 ;
        RECT 1.1910 0.0300 1.2410 0.3820 ;
        RECT 1.4950 0.0300 1.5450 0.5660 ;
        RECT 1.7990 0.0300 1.8490 0.3820 ;
        RECT 0.8870 0.0300 0.9370 0.3820 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 7.2960 3.3740 ;
    END
  END VSS

  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7950 0.6560 1.4850 0.7160 ;
        RECT 0.9740 0.7160 1.1340 0.8150 ;
    END
    ANTENNAGATEAREA 0.183 ;
  END SLEEP

  PIN SLEEPOUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9510 1.1400 2.0010 1.3580 ;
        RECT 1.6470 1.1400 1.6970 1.3580 ;
        RECT 1.6470 1.0800 2.0010 1.1400 ;
        RECT 1.6470 1.0730 1.6970 1.0800 ;
        RECT 4.0790 0.8660 4.1290 1.3580 ;
        RECT 6.2070 0.8660 6.2570 1.3580 ;
        RECT 5.9030 0.8660 5.9530 1.3580 ;
        RECT 5.5990 0.8660 5.6490 1.3580 ;
        RECT 5.2950 0.8660 5.3450 1.3580 ;
        RECT 4.9910 0.8660 5.0410 1.3580 ;
        RECT 4.6870 0.8660 4.7370 1.3580 ;
        RECT 4.3830 0.8660 4.4330 1.3580 ;
        RECT 2.2550 0.8660 2.3050 1.3580 ;
        RECT 2.5590 0.8660 2.6090 1.3580 ;
        RECT 2.8630 0.8660 2.9130 1.3580 ;
        RECT 3.1670 0.8660 3.2170 1.3580 ;
        RECT 3.4710 0.8660 3.5210 1.3580 ;
        RECT 3.7750 0.8660 3.8250 1.3580 ;
        RECT 1.9510 0.8660 2.0010 1.0800 ;
        RECT 1.9510 0.8060 6.5270 0.8660 ;
        RECT 4.0790 0.7950 4.1290 0.8060 ;
        RECT 6.2070 0.7950 6.2570 0.8060 ;
        RECT 5.9030 0.7950 5.9530 0.8060 ;
        RECT 5.5990 0.7950 5.6490 0.8060 ;
        RECT 5.2950 0.7950 5.3450 0.8060 ;
        RECT 4.9910 0.7950 5.0410 0.8060 ;
        RECT 4.6870 0.7950 4.7370 0.8060 ;
        RECT 4.3830 0.7950 4.4330 0.8060 ;
        RECT 1.9510 0.7950 2.0010 0.8060 ;
        RECT 2.2550 0.7950 2.3050 0.8060 ;
        RECT 2.5590 0.7950 2.6090 0.8060 ;
        RECT 2.8630 0.7950 2.9130 0.8060 ;
        RECT 3.1670 0.7950 3.2170 0.8060 ;
        RECT 3.4710 0.7950 3.5210 0.8060 ;
        RECT 3.7750 0.7950 3.8250 0.8060 ;
        RECT 6.4770 0.6630 6.5270 0.8060 ;
        RECT 6.4700 0.5620 6.5930 0.6630 ;
        RECT 1.6470 0.5520 6.5930 0.5620 ;
        RECT 1.6470 0.5020 6.5870 0.5520 ;
        RECT 4.0790 0.1790 4.1290 0.5020 ;
        RECT 4.6870 0.1790 4.7370 0.5020 ;
        RECT 4.9910 0.1790 5.0410 0.5020 ;
        RECT 5.2950 0.1790 5.3450 0.5020 ;
        RECT 5.5990 0.1790 5.6490 0.5020 ;
        RECT 5.9030 0.1790 5.9530 0.5020 ;
        RECT 6.2070 0.1790 6.2570 0.5020 ;
        RECT 4.3830 0.1790 4.4330 0.5020 ;
        RECT 1.6470 0.1800 1.6970 0.5020 ;
        RECT 1.9510 0.1800 2.0010 0.5020 ;
        RECT 2.2550 0.1800 2.3050 0.5020 ;
        RECT 2.5590 0.1790 2.6090 0.5020 ;
        RECT 2.8630 0.1790 2.9130 0.5020 ;
        RECT 3.1670 0.1790 3.2170 0.5020 ;
        RECT 3.4710 0.1790 3.5210 0.5020 ;
        RECT 3.7750 0.1790 3.8250 0.5020 ;
    END
    ANTENNADIFFAREA 2.3808 ;
  END SLEEPOUT

  PIN VDDG
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 6.2900 2.0730 6.4800 2.1830 ;
        RECT 6.3560 2.0110 6.4160 2.0730 ;
        RECT 6.3560 2.1830 6.4160 2.4930 ;
        RECT 1.3420 2.4930 6.6530 2.5430 ;
        RECT 3.4710 1.8370 3.5210 2.4930 ;
        RECT 3.1670 1.8370 3.2170 2.4930 ;
        RECT 2.8630 1.8370 2.9130 2.4930 ;
        RECT 2.5590 1.8370 2.6090 2.4930 ;
        RECT 2.2550 1.8370 2.3050 2.4930 ;
        RECT 1.9510 1.8370 2.0010 2.4930 ;
        RECT 1.6470 1.8370 1.6970 2.4930 ;
        RECT 1.3430 1.8370 1.3930 2.4930 ;
        RECT 3.7750 1.8370 3.8250 2.4930 ;
        RECT 4.0790 1.8370 4.1290 2.4930 ;
        RECT 4.3830 1.8370 4.4330 2.4930 ;
        RECT 4.6870 1.8370 4.7370 2.4930 ;
        RECT 4.9910 1.8370 5.0410 2.4930 ;
        RECT 5.2950 1.8370 5.3450 2.4930 ;
        RECT 5.5990 1.8370 5.6490 2.4930 ;
        RECT 5.9030 1.8370 5.9530 2.4930 ;
    END
  END VDDG

  PIN VDD
    DIRECTION OUTPUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 7.2960 1.7020 ;
        RECT 3.6230 1.7020 3.6730 2.3090 ;
        RECT 3.3190 1.7020 3.3690 2.3090 ;
        RECT 3.0150 1.7020 3.0650 2.3090 ;
        RECT 2.7110 1.7020 2.7610 2.3100 ;
        RECT 2.4070 1.7020 2.4570 2.3100 ;
        RECT 2.1030 1.7020 2.1530 2.3100 ;
        RECT 1.7990 1.7020 1.8490 2.3100 ;
        RECT 1.1910 1.7020 1.2410 2.4940 ;
        RECT 1.4950 1.7020 1.5450 2.3100 ;
        RECT 3.9270 1.7020 3.9770 2.3100 ;
        RECT 4.2310 1.7020 4.2810 2.3100 ;
        RECT 4.5350 1.7020 4.5850 2.3100 ;
        RECT 4.8390 1.7020 4.8890 2.3100 ;
        RECT 5.1430 1.7020 5.1930 2.3100 ;
        RECT 5.4470 1.7020 5.4970 2.3090 ;
        RECT 5.7510 1.7020 5.8010 2.3090 ;
        RECT 6.0550 1.7020 6.1050 2.3090 ;
    END
  END VDD
  OBS
    LAYER PO ;
      RECT 1.7330 1.7070 1.7630 3.2330 ;
      RECT 1.1250 1.7070 1.1550 3.2330 ;
      RECT 1.1250 0.1190 1.1550 1.6070 ;
      RECT 1.4290 1.7070 1.4590 3.2330 ;
      RECT 1.8850 0.1200 1.9150 1.6070 ;
      RECT 3.8610 1.7070 3.8910 3.2330 ;
      RECT 1.2770 0.1200 1.3070 1.6070 ;
      RECT 1.7330 0.1200 1.7630 1.6070 ;
      RECT 0.9730 1.7070 1.0030 3.2330 ;
      RECT 1.4290 0.1200 1.4590 1.6070 ;
      RECT 1.5810 0.1200 1.6110 1.6070 ;
      RECT 1.5810 1.7070 1.6110 3.2330 ;
      RECT 7.2050 0.1200 7.2350 1.6070 ;
      RECT 6.9010 0.1200 6.9310 1.6070 ;
      RECT 6.7490 0.1200 6.7790 1.6070 ;
      RECT 7.0530 0.1200 7.0830 1.6070 ;
      RECT 6.7490 1.7070 6.7790 3.2290 ;
      RECT 6.9010 1.7070 6.9310 3.2290 ;
      RECT 7.0530 1.7070 7.0830 3.2290 ;
      RECT 7.2050 1.7070 7.2350 3.2290 ;
      RECT 0.3650 0.1190 0.3950 1.6070 ;
      RECT 0.0610 0.1200 0.0910 1.6070 ;
      RECT 0.2130 0.1200 0.2430 1.6070 ;
      RECT 0.5170 0.1200 0.5470 1.6070 ;
      RECT 0.0610 1.7070 0.0910 3.2330 ;
      RECT 0.5170 1.7070 0.5470 3.2330 ;
      RECT 0.3650 1.7070 0.3950 3.2330 ;
      RECT 0.2130 1.7070 0.2430 3.2330 ;
      RECT 4.1650 1.7070 4.1950 3.2330 ;
      RECT 4.3170 1.7070 4.3470 3.2330 ;
      RECT 4.4690 1.7070 4.4990 3.2330 ;
      RECT 4.6210 1.7070 4.6510 3.2330 ;
      RECT 4.7730 1.7070 4.8030 3.2330 ;
      RECT 4.9250 1.7070 4.9550 3.2330 ;
      RECT 5.0770 1.7070 5.1070 3.2330 ;
      RECT 5.2290 1.7070 5.2590 3.2330 ;
      RECT 5.3810 1.7070 5.4110 3.2330 ;
      RECT 5.5330 1.7070 5.5630 3.2290 ;
      RECT 5.6850 1.7070 5.7150 3.2290 ;
      RECT 5.8370 1.7070 5.8670 3.2290 ;
      RECT 5.9890 1.7070 6.0190 3.2290 ;
      RECT 6.1410 1.7070 6.1710 3.2290 ;
      RECT 6.2930 1.7070 6.3230 3.2290 ;
      RECT 6.4450 1.7070 6.4750 3.2290 ;
      RECT 4.1650 0.1200 4.1950 1.6070 ;
      RECT 4.3170 0.1200 4.3470 1.6070 ;
      RECT 4.4690 0.1200 4.4990 1.6070 ;
      RECT 4.6210 0.1200 4.6510 1.6070 ;
      RECT 4.7730 0.1200 4.8030 1.6070 ;
      RECT 4.9250 0.1200 4.9550 1.6070 ;
      RECT 5.0770 0.1200 5.1070 1.6070 ;
      RECT 5.2290 0.1200 5.2590 1.6070 ;
      RECT 5.3810 0.1200 5.4110 1.6070 ;
      RECT 5.5330 0.1200 5.5630 1.6070 ;
      RECT 6.4450 0.1200 6.4750 1.6070 ;
      RECT 6.1410 0.1200 6.1710 1.6070 ;
      RECT 5.9890 0.1200 6.0190 1.6070 ;
      RECT 5.8370 0.1200 5.8670 1.6070 ;
      RECT 5.6850 0.1200 5.7150 1.6070 ;
      RECT 2.6450 1.7070 2.6750 3.2290 ;
      RECT 2.7970 1.7070 2.8270 3.2290 ;
      RECT 2.9490 1.7070 2.9790 3.2290 ;
      RECT 3.1010 1.7070 3.1310 3.2290 ;
      RECT 3.2530 1.7070 3.2830 3.2290 ;
      RECT 3.4050 1.7070 3.4350 3.2290 ;
      RECT 3.5570 1.7070 3.5870 3.2290 ;
      RECT 3.7090 1.7070 3.7390 3.2290 ;
      RECT 3.4050 0.1200 3.4350 1.6070 ;
      RECT 3.2530 0.1200 3.2830 1.6070 ;
      RECT 3.1010 0.1200 3.1310 1.6070 ;
      RECT 2.9490 0.1200 2.9790 1.6070 ;
      RECT 3.5570 0.1200 3.5870 1.6070 ;
      RECT 3.7090 0.1200 3.7390 1.6070 ;
      RECT 3.8610 0.1200 3.8910 1.6070 ;
      RECT 4.0130 0.1200 4.0430 1.6070 ;
      RECT 6.2930 0.1200 6.3230 1.6070 ;
      RECT 4.0130 1.7070 4.0430 3.2330 ;
      RECT 2.7970 0.1200 2.8270 1.6070 ;
      RECT 2.4930 0.1200 2.5230 1.6070 ;
      RECT 2.1890 1.7070 2.2190 3.2330 ;
      RECT 2.1890 0.1200 2.2190 1.6070 ;
      RECT 2.6450 0.1200 2.6750 1.6070 ;
      RECT 2.0370 0.1200 2.0670 1.6070 ;
      RECT 2.3410 1.7070 2.3710 3.2330 ;
      RECT 2.4930 1.7070 2.5230 3.2330 ;
      RECT 0.6690 0.1200 0.6990 3.2330 ;
      RECT 6.5970 0.1200 6.6270 3.2330 ;
      RECT 0.8210 0.1200 0.8510 1.6070 ;
      RECT 2.3410 0.1200 2.3710 1.6070 ;
      RECT 0.8210 1.7070 0.8510 3.2330 ;
      RECT 2.0370 1.7070 2.0670 3.2330 ;
      RECT 0.9730 0.1200 1.0030 1.6070 ;
      RECT 1.2770 1.7070 1.3070 3.2330 ;
      RECT 1.8850 1.7070 1.9150 3.2330 ;
    LAYER NWELL ;
      RECT 0.5710 0.6790 6.7170 2.6650 ;
    LAYER M1 ;
      RECT 0.8870 1.4590 6.6530 1.5190 ;
      RECT 6.3590 1.0480 6.4090 1.4590 ;
      RECT 1.4950 1.0480 1.5450 1.4590 ;
      RECT 0.8870 1.0480 0.9370 1.4590 ;
      RECT 1.1910 1.0480 1.2410 1.4590 ;
      RECT 1.7990 1.2340 1.8490 1.4590 ;
      RECT 2.1030 1.0480 2.1530 1.4590 ;
      RECT 2.4070 1.0480 2.4570 1.4590 ;
      RECT 2.7110 1.0480 2.7610 1.4590 ;
      RECT 3.0150 1.0480 3.0650 1.4590 ;
      RECT 3.3190 1.0480 3.3690 1.4590 ;
      RECT 3.6230 1.0480 3.6730 1.4590 ;
      RECT 3.9270 1.0480 3.9770 1.4590 ;
      RECT 4.2310 1.0480 4.2810 1.4590 ;
      RECT 4.5350 1.0480 4.5850 1.4590 ;
      RECT 4.8390 1.0480 4.8890 1.4590 ;
      RECT 5.1430 1.0480 5.1930 1.4590 ;
      RECT 5.4470 1.0480 5.4970 1.4590 ;
      RECT 5.7510 1.0480 5.8010 1.4590 ;
      RECT 6.0550 1.0480 6.1050 1.4590 ;
      RECT 1.5550 0.6560 6.3490 0.7160 ;
      RECT 1.0390 0.9600 1.0890 1.3580 ;
      RECT 1.0390 0.1800 1.0890 0.5020 ;
      RECT 1.3430 0.9600 1.3930 1.3580 ;
      RECT 1.3430 0.7950 1.3930 0.9000 ;
      RECT 0.6590 0.5020 1.3930 0.5620 ;
      RECT 1.3430 0.1800 1.3930 0.5020 ;
      RECT 1.5710 0.7160 1.6210 0.9000 ;
      RECT 0.6590 0.9000 1.6210 0.9600 ;
      RECT 0.6590 0.5620 0.7090 0.9000 ;
      RECT 0.7350 0.9600 0.7850 1.3580 ;
      RECT 0.7350 0.1800 0.7850 0.5020 ;
      RECT 0.6430 2.6030 6.0450 2.6530 ;
  END
END HEAD2X32_LVT

MACRO HEAD2X4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.584 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SLEEPOUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1910 1.0840 1.5450 1.1440 ;
        RECT 1.1910 1.1440 1.2410 1.4030 ;
        RECT 1.4950 1.1440 1.5450 1.3580 ;
        RECT 1.4950 0.8660 1.5450 1.0840 ;
        RECT 1.4950 0.8060 1.8040 0.8660 ;
        RECT 1.4950 0.7950 1.5450 0.8060 ;
        RECT 1.7540 0.6630 1.8040 0.8060 ;
        RECT 1.7540 0.5620 1.8790 0.6630 ;
        RECT 1.1910 0.5520 1.8790 0.5620 ;
        RECT 1.1910 0.5020 1.8750 0.5520 ;
        RECT 1.1910 0.1800 1.2410 0.5020 ;
        RECT 1.4950 0.1800 1.5450 0.5020 ;
    END
    ANTENNADIFFAREA 0.2976 ;
  END SLEEPOUT

  PIN VDDG
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 1.5760 2.0730 1.7660 2.1830 ;
        RECT 1.6420 2.0110 1.7020 2.0730 ;
        RECT 1.6420 2.1830 1.7020 2.4930 ;
        RECT 0.8860 2.4930 1.9410 2.5430 ;
        RECT 1.1910 1.8370 1.2410 2.4930 ;
        RECT 0.8870 1.8370 0.9370 2.4930 ;
    END
  END VDDG

  PIN VDD
    DIRECTION OUTPUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.5840 1.7020 ;
        RECT 1.3430 1.7020 1.3930 2.3100 ;
        RECT 0.7350 1.7020 0.7850 2.4940 ;
        RECT 1.0390 1.7020 1.0890 2.3100 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.5840 0.0300 ;
        RECT 1.6470 0.0300 1.6970 0.3820 ;
        RECT 1.0390 0.0300 1.0890 0.5660 ;
        RECT 1.3430 0.0300 1.3930 0.3820 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 2.5840 3.3740 ;
    END
  END VSS

  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8530 0.6450 1.0280 0.8150 ;
    END
    ANTENNAGATEAREA 0.0366 ;
  END SLEEP
  OBS
    LAYER NWELL ;
      RECT 0.5710 0.6790 1.9760 2.6650 ;
    LAYER M1 ;
      RECT 1.0390 1.4590 1.9410 1.5190 ;
      RECT 1.6470 1.0480 1.6970 1.4590 ;
      RECT 1.0390 1.1400 1.0890 1.4590 ;
      RECT 1.3430 1.2340 1.3930 1.4590 ;
      RECT 1.0990 0.6560 1.6370 0.7160 ;
      RECT 0.8870 1.0210 0.9370 1.5040 ;
      RECT 0.8870 0.9600 0.9370 0.9610 ;
      RECT 0.6590 0.5020 0.9370 0.5620 ;
      RECT 0.8870 0.1800 0.9370 0.5020 ;
      RECT 1.1150 0.7160 1.1650 0.9610 ;
      RECT 0.6590 0.9610 1.1650 1.0210 ;
      RECT 0.6590 0.5620 0.7090 0.9610 ;
      RECT 0.6430 2.6030 1.3330 2.6530 ;
    LAYER PO ;
      RECT 2.4930 1.7160 2.5230 3.2300 ;
      RECT 2.4930 0.1200 2.5230 1.6070 ;
      RECT 2.3410 0.1200 2.3710 1.6070 ;
      RECT 2.1890 0.1200 2.2190 1.6070 ;
      RECT 2.0370 0.1200 2.0670 1.6070 ;
      RECT 0.0610 0.1200 0.0910 1.6070 ;
      RECT 0.5170 0.1200 0.5470 1.6070 ;
      RECT 0.2130 0.1200 0.2430 1.6070 ;
      RECT 0.3650 0.1200 0.3950 1.6070 ;
      RECT 2.3410 1.7210 2.3710 3.2310 ;
      RECT 2.1890 1.7210 2.2190 3.2310 ;
      RECT 2.0370 1.7210 2.0670 3.2310 ;
      RECT 0.0610 1.7070 0.0910 3.2350 ;
      RECT 0.2130 1.7070 0.2430 3.2350 ;
      RECT 0.3650 1.7070 0.3950 3.2350 ;
      RECT 0.5170 1.7070 0.5470 3.2350 ;
      RECT 1.7330 1.7070 1.7630 3.2310 ;
      RECT 1.7330 0.1200 1.7630 1.6070 ;
      RECT 1.5810 0.1200 1.6110 1.6070 ;
      RECT 1.8850 0.1200 1.9150 3.2310 ;
      RECT 1.5810 1.7210 1.6110 3.2310 ;
      RECT 0.8210 1.7070 0.8510 3.2350 ;
      RECT 1.4290 1.7210 1.4590 3.2310 ;
      RECT 1.2770 1.7070 1.3070 3.2350 ;
      RECT 0.6690 0.1190 0.6990 3.2350 ;
      RECT 0.9730 1.7070 1.0030 3.2350 ;
      RECT 1.4290 0.1200 1.4590 1.6070 ;
      RECT 0.8210 0.1200 0.8510 1.6070 ;
      RECT 1.2770 0.1200 1.3070 1.6070 ;
      RECT 0.9730 0.1200 1.0030 1.6070 ;
      RECT 1.1250 0.1200 1.1550 1.6070 ;
      RECT 1.1250 1.7070 1.1550 3.2350 ;
  END
END HEAD2X4_LVT

MACRO HEAD2X8_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.192 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SLEEPOUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1910 0.5020 2.4830 0.5520 ;
        RECT 1.1910 0.1800 1.2410 0.5020 ;
        RECT 1.1910 0.5520 2.4890 0.5620 ;
        RECT 2.1030 0.1790 2.1530 0.5020 ;
        RECT 1.7990 0.1800 1.8490 0.5020 ;
        RECT 1.4950 0.1800 1.5450 0.5020 ;
        RECT 2.3650 0.5620 2.4890 0.6630 ;
        RECT 2.3650 0.6630 2.4150 0.8060 ;
        RECT 1.4950 0.8060 2.4150 0.8660 ;
        RECT 2.1030 0.8660 2.1530 1.3580 ;
        RECT 2.1030 0.7950 2.1530 0.8060 ;
        RECT 1.7990 0.8660 1.8490 1.3580 ;
        RECT 1.7990 0.7950 1.8490 0.8060 ;
        RECT 1.4950 0.7950 1.5450 0.8060 ;
        RECT 1.4950 0.8660 1.5450 1.0840 ;
        RECT 1.1910 1.0840 1.5450 1.1440 ;
        RECT 1.1910 1.1440 1.2410 1.3580 ;
        RECT 1.1910 1.0730 1.2410 1.0840 ;
        RECT 1.4950 1.1440 1.5450 1.3580 ;
    END
    ANTENNADIFFAREA 0.5952 ;
  END SLEEPOUT

  PIN VDDG
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 2.1840 2.0730 2.3740 2.1830 ;
        RECT 2.2500 2.0110 2.3100 2.0730 ;
        RECT 2.2500 2.1830 2.3100 2.4930 ;
        RECT 0.8860 2.4930 2.5490 2.5430 ;
        RECT 0.8870 1.8370 0.9370 2.4930 ;
        RECT 1.7990 1.8370 1.8490 2.4930 ;
        RECT 1.4950 1.8370 1.5450 2.4930 ;
        RECT 1.1910 1.8370 1.2410 2.4930 ;
    END
  END VDDG

  PIN VDD
    DIRECTION OUTPUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.1920 1.7020 ;
        RECT 0.7350 1.7020 0.7850 2.4940 ;
        RECT 1.0390 1.7020 1.0890 2.3100 ;
        RECT 1.9510 1.7020 2.0010 2.3100 ;
        RECT 1.6470 1.7020 1.6970 2.3100 ;
        RECT 1.3430 1.7020 1.3930 2.3100 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.1920 0.0300 ;
        RECT 1.0390 0.0300 1.0890 0.5660 ;
        RECT 1.3430 0.0300 1.3930 0.3820 ;
        RECT 0.7350 0.0300 0.7850 0.3790 ;
        RECT 2.2550 0.0300 2.3050 0.3820 ;
        RECT 1.9510 0.0300 2.0010 0.3820 ;
        RECT 1.6470 0.0300 1.6970 0.3820 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 3.1920 3.3740 ;
    END
  END VSS

  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7950 0.6560 1.0290 0.7160 ;
        RECT 0.8340 0.7160 0.9940 0.8150 ;
    END
    ANTENNAGATEAREA 0.0732 ;
  END SLEEP
  OBS
    LAYER NWELL ;
      RECT 0.5710 0.6790 2.5840 2.6650 ;
    LAYER M1 ;
      RECT 0.7350 1.4590 2.5490 1.5190 ;
      RECT 2.2550 1.0480 2.3050 1.4590 ;
      RECT 1.0390 1.0980 1.0890 1.4590 ;
      RECT 0.7350 1.0980 0.7850 1.4590 ;
      RECT 1.3430 1.2340 1.3930 1.4590 ;
      RECT 1.6470 1.0480 1.6970 1.4590 ;
      RECT 1.9510 1.0480 2.0010 1.4590 ;
      RECT 1.0990 0.6560 2.2450 0.7160 ;
      RECT 0.8870 0.9890 0.9370 1.3270 ;
      RECT 0.8870 0.8730 0.9370 0.9290 ;
      RECT 0.5070 0.5320 0.9370 0.5620 ;
      RECT 0.5080 0.5020 0.9370 0.5320 ;
      RECT 0.8870 0.1800 0.9370 0.5020 ;
      RECT 1.1150 0.7160 1.1650 0.9290 ;
      RECT 0.5070 0.9290 1.1650 0.9890 ;
      RECT 0.5070 0.5620 0.5570 0.9290 ;
      RECT 0.4910 2.6030 1.9410 2.6530 ;
    LAYER PO ;
      RECT 0.0610 0.1200 0.0910 1.6070 ;
      RECT 0.2130 0.1200 0.2430 1.6070 ;
      RECT 0.3650 0.1200 0.3950 1.6070 ;
      RECT 3.1010 0.1200 3.1310 1.6070 ;
      RECT 2.7970 0.1200 2.8270 1.6070 ;
      RECT 2.9490 0.1200 2.9790 1.6070 ;
      RECT 2.6450 0.1200 2.6750 1.6070 ;
      RECT 3.1010 1.7070 3.1310 3.2350 ;
      RECT 2.7970 1.7070 2.8270 3.2350 ;
      RECT 2.6450 1.7070 2.6750 3.2350 ;
      RECT 2.9490 1.7070 2.9790 3.2350 ;
      RECT 0.2130 1.7070 0.2430 3.2350 ;
      RECT 0.0610 1.7070 0.0910 3.2350 ;
      RECT 0.3650 1.7070 0.3950 3.2350 ;
      RECT 2.3410 1.7070 2.3710 3.2340 ;
      RECT 2.3410 0.1200 2.3710 1.6070 ;
      RECT 2.0370 0.1200 2.0670 1.6070 ;
      RECT 1.7330 1.7070 1.7630 3.2350 ;
      RECT 1.7330 0.1200 1.7630 1.6070 ;
      RECT 2.1890 0.1200 2.2190 1.6070 ;
      RECT 1.5810 0.1200 1.6110 1.6070 ;
      RECT 1.8850 1.7070 1.9150 3.2350 ;
      RECT 2.0370 1.7070 2.0670 3.2340 ;
      RECT 2.4930 0.1200 2.5230 3.2340 ;
      RECT 1.8850 0.1200 1.9150 1.6070 ;
      RECT 1.5810 1.7070 1.6110 3.2350 ;
      RECT 0.5170 0.1200 0.5470 3.2350 ;
      RECT 0.8210 1.7070 0.8510 3.2350 ;
      RECT 1.4290 1.7070 1.4590 3.2350 ;
      RECT 1.2770 1.7070 1.3070 3.2350 ;
      RECT 0.6690 1.7070 0.6990 3.2350 ;
      RECT 0.6690 0.1200 0.6990 1.6070 ;
      RECT 0.9730 1.7070 1.0030 3.2350 ;
      RECT 1.4290 0.1200 1.4590 1.6070 ;
      RECT 2.1890 1.7070 2.2190 3.2340 ;
      RECT 0.8210 0.1200 0.8510 1.6070 ;
      RECT 1.2770 0.1200 1.3070 1.6070 ;
      RECT 0.9730 0.1200 1.0030 1.6070 ;
      RECT 1.1250 0.1200 1.1550 1.6070 ;
      RECT 1.1250 1.7070 1.1550 3.2350 ;
  END
END HEAD2X8_LVT

MACRO HEADX16_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.256 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDDG
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.6660 1.0090 0.8560 1.1190 ;
        RECT 0.7300 1.1190 0.7900 1.1650 ;
        RECT 0.7300 0.8810 0.7900 1.0090 ;
        RECT 0.7300 0.8450 3.3690 0.8810 ;
        RECT 0.7350 0.8310 3.3690 0.8450 ;
        RECT 1.7990 0.8810 1.8490 1.5610 ;
        RECT 1.4950 0.8810 1.5450 1.5610 ;
        RECT 1.1910 0.8810 1.2410 1.5610 ;
        RECT 2.1030 0.8810 2.1530 1.5610 ;
        RECT 2.4070 0.8810 2.4570 1.5610 ;
        RECT 2.7110 0.8810 2.7610 1.5610 ;
        RECT 3.0150 0.8810 3.0650 1.5610 ;
        RECT 3.3190 0.8810 3.3690 1.5610 ;
    END
  END VDDG

  PIN VDD
    DIRECTION OUTPUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.2560 1.7020 ;
        RECT 1.3430 1.0150 1.3930 1.6420 ;
        RECT 3.4710 0.8310 3.5210 1.6420 ;
        RECT 3.1670 1.0150 3.2170 1.6420 ;
        RECT 2.8630 1.0150 2.9130 1.6420 ;
        RECT 2.5590 1.0150 2.6090 1.6420 ;
        RECT 2.2550 1.0150 2.3050 1.6420 ;
        RECT 1.9510 1.0150 2.0010 1.6420 ;
        RECT 1.0390 1.0150 1.0890 1.6420 ;
        RECT 1.6470 1.0150 1.6970 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.2560 0.0300 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 4.2560 3.3740 ;
    END
  END VSS

  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0990 0.6700 3.4610 0.7300 ;
        RECT 1.1200 0.5530 1.3100 0.6700 ;
    END
  END SLEEP
  OBS
    LAYER NWELL ;
      RECT 0.5710 0.6790 3.6770 2.6650 ;
    LAYER PO ;
      RECT 4.1650 0.1230 4.1950 1.6210 ;
      RECT 3.7090 0.1230 3.7390 1.6210 ;
      RECT 3.8610 0.1230 3.8910 1.6210 ;
      RECT 4.0130 0.1230 4.0430 1.6210 ;
      RECT 0.5170 0.1230 0.5470 1.6210 ;
      RECT 0.3650 0.1230 0.3950 1.6210 ;
      RECT 0.2130 0.1230 0.2430 1.6210 ;
      RECT 0.0610 0.1230 0.0910 1.6210 ;
      RECT 0.0610 1.7240 0.0910 3.2220 ;
      RECT 0.5170 1.7230 0.5470 3.2210 ;
      RECT 0.3650 1.7230 0.3950 3.2210 ;
      RECT 0.2130 1.7230 0.2430 3.2210 ;
      RECT 4.1650 1.7230 4.1950 3.2210 ;
      RECT 3.7090 1.7230 3.7390 3.2210 ;
      RECT 3.8610 1.7230 3.8910 3.2210 ;
      RECT 4.0130 1.7230 4.0430 3.2210 ;
      RECT 1.2770 1.7230 1.3070 3.2210 ;
      RECT 1.1250 1.7230 1.1550 3.2210 ;
      RECT 1.7330 1.7230 1.7630 3.2210 ;
      RECT 1.4290 1.7230 1.4590 3.2210 ;
      RECT 0.9730 1.7230 1.0030 3.2210 ;
      RECT 0.8210 1.7230 0.8510 3.2210 ;
      RECT 1.5810 1.7230 1.6110 3.2210 ;
      RECT 0.6690 1.7240 0.6990 3.2220 ;
      RECT 1.8850 1.7230 1.9150 3.2210 ;
      RECT 2.0370 1.7230 2.0670 3.2210 ;
      RECT 2.1890 1.7230 2.2190 3.2210 ;
      RECT 2.3410 1.7230 2.3710 3.2210 ;
      RECT 3.5570 1.7230 3.5870 3.2210 ;
      RECT 2.4930 1.7230 2.5230 3.2210 ;
      RECT 2.6450 1.7230 2.6750 3.2210 ;
      RECT 2.7970 1.7230 2.8270 3.2210 ;
      RECT 2.9490 1.7230 2.9790 3.2210 ;
      RECT 3.1010 1.7230 3.1310 3.2210 ;
      RECT 3.2530 1.7230 3.2830 3.2210 ;
      RECT 3.4050 1.7230 3.4350 3.2210 ;
      RECT 3.4050 0.1230 3.4350 1.6210 ;
      RECT 3.2530 0.1230 3.2830 1.6210 ;
      RECT 3.1010 0.1230 3.1310 1.6210 ;
      RECT 2.9490 0.1230 2.9790 1.6210 ;
      RECT 2.7970 0.1230 2.8270 1.6210 ;
      RECT 2.6450 0.1230 2.6750 1.6210 ;
      RECT 2.4930 0.1230 2.5230 1.6210 ;
      RECT 3.5570 0.1230 3.5870 1.6210 ;
      RECT 2.3410 0.1230 2.3710 1.6210 ;
      RECT 2.1890 0.1230 2.2190 1.6210 ;
      RECT 2.0370 0.1230 2.0670 1.6210 ;
      RECT 1.8850 0.1230 1.9150 1.6210 ;
      RECT 0.6690 0.1230 0.6990 1.6210 ;
      RECT 1.5810 0.1230 1.6110 1.6210 ;
      RECT 0.8210 0.1230 0.8510 1.6210 ;
      RECT 0.9730 0.1230 1.0030 1.6210 ;
      RECT 1.4290 0.1230 1.4590 1.6210 ;
      RECT 1.7330 0.1230 1.7630 1.6210 ;
      RECT 1.1250 0.1230 1.1550 1.6210 ;
      RECT 1.2770 0.1230 1.3070 1.6210 ;
  END
END HEADX16_LVT

MACRO DFFSSRX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.712 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.5050 0.2170 4.6150 0.2700 ;
        RECT 4.2310 0.2700 4.6150 0.3200 ;
        RECT 4.5050 0.3200 4.6150 0.3590 ;
        RECT 4.2310 0.1480 4.2810 0.2700 ;
        RECT 4.5470 0.3590 4.5970 0.9180 ;
        RECT 4.2310 0.9180 4.5970 0.9680 ;
        RECT 4.2310 0.9680 4.2810 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.9270 0.1480 3.9770 0.3940 ;
        RECT 3.9270 0.3940 4.4350 0.4010 ;
        RECT 3.9270 0.4010 4.4730 0.4440 ;
        RECT 4.3530 0.4440 4.4730 0.5110 ;
        RECT 4.4230 0.5110 4.4730 0.8040 ;
        RECT 3.9270 0.8040 4.4730 0.8540 ;
        RECT 3.9270 0.8540 3.9770 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.7120 1.7020 ;
        RECT 3.7750 0.9120 3.8250 1.6420 ;
        RECT 4.0790 0.9600 4.1290 1.6420 ;
        RECT 4.3830 1.0520 4.4330 1.6420 ;
        RECT 3.6630 1.4660 3.7130 1.6420 ;
        RECT 0.2790 1.3460 0.3290 1.6420 ;
        RECT 1.4050 1.3660 1.4550 1.6420 ;
        RECT 2.4070 1.3660 2.4570 1.6420 ;
        RECT 3.1510 1.4160 3.7130 1.4660 ;
        RECT 0.2790 1.2960 0.6330 1.3460 ;
        RECT 1.3050 1.3160 1.4550 1.3660 ;
        RECT 2.2550 1.3160 2.4570 1.3660 ;
        RECT 3.6230 1.1920 3.6730 1.4160 ;
        RECT 0.2790 0.9300 0.3290 1.2960 ;
        RECT 0.5830 0.9800 0.6330 1.2960 ;
        RECT 2.2550 1.1000 2.3050 1.3160 ;
    END
  END VDD

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7010 0.4210 0.7510 ;
        RECT 0.2490 0.7510 0.3590 0.8250 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SETB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.4650 1.3330 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.7120 0.0300 ;
        RECT 3.1270 0.0300 3.1770 0.2040 ;
        RECT 0.2790 0.0300 0.3290 0.3550 ;
        RECT 3.6230 0.0300 3.6730 0.4010 ;
        RECT 3.7750 0.0300 3.8250 0.4080 ;
        RECT 4.0790 0.0300 4.1290 0.3190 ;
        RECT 4.3830 0.0300 4.4330 0.2200 ;
        RECT 2.0270 0.0300 2.0770 0.3010 ;
        RECT 3.1270 0.2040 3.2330 0.2540 ;
        RECT 0.2790 0.3550 0.6330 0.4050 ;
        RECT 1.3430 0.3010 2.4570 0.3510 ;
        RECT 0.5830 0.4050 0.6330 0.5290 ;
        RECT 0.2790 0.4050 0.3290 0.5130 ;
        RECT 2.4070 0.3510 2.4570 0.4750 ;
        RECT 1.3430 0.3510 1.3930 0.5760 ;
        RECT 2.2550 0.3510 2.3050 0.4750 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9470 0.8670 1.1190 0.9770 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 0.1070 0.5110 0.2010 ;
        RECT 0.4010 0.2010 0.7250 0.2510 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END RSTB
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 4.8270 1.7730 ;
    LAYER M1 ;
      RECT 0.4310 0.8440 0.7500 0.8940 ;
      RECT 0.7000 0.6230 0.7500 0.8440 ;
      RECT 0.7000 0.5730 0.8770 0.6230 ;
      RECT 0.4310 0.4550 0.4810 0.6010 ;
      RECT 0.4310 0.8940 0.4810 1.2460 ;
      RECT 0.4310 0.6010 0.5210 0.6510 ;
      RECT 0.4710 0.6510 0.5210 0.8440 ;
      RECT 2.9230 1.5280 3.6130 1.5780 ;
      RECT 4.1360 0.6540 4.1860 0.7040 ;
      RECT 4.1360 0.6040 4.3730 0.6540 ;
      RECT 3.6800 0.7040 4.1860 0.7540 ;
      RECT 3.3790 0.5770 3.7300 0.6270 ;
      RECT 3.6800 0.6270 3.7300 0.7040 ;
      RECT 3.6800 0.7540 3.7300 0.7580 ;
      RECT 0.7190 0.3010 1.1050 0.3510 ;
      RECT 0.7350 1.3160 1.1060 1.3660 ;
      RECT 0.7350 0.9800 0.7850 1.3160 ;
      RECT 1.0990 0.1040 1.9410 0.1540 ;
      RECT 1.7230 0.1540 1.7730 0.2170 ;
      RECT 1.8590 1.4170 2.2450 1.4670 ;
      RECT 1.4950 0.7260 1.5970 0.7760 ;
      RECT 1.4950 0.7760 1.5450 1.1520 ;
      RECT 1.5470 0.6760 1.5970 0.7260 ;
      RECT 1.5470 0.6260 1.6370 0.6760 ;
      RECT 1.5470 0.4960 1.5970 0.6260 ;
      RECT 1.4790 0.4460 1.5970 0.4960 ;
      RECT 3.8120 0.6040 4.0690 0.6540 ;
      RECT 2.8630 0.3000 2.9130 1.2160 ;
      RECT 3.2790 0.5270 3.3290 0.6540 ;
      RECT 3.0750 0.6540 3.3290 0.6770 ;
      RECT 3.0750 0.6770 3.4090 0.7040 ;
      RECT 3.2790 0.7040 3.4090 0.7270 ;
      RECT 3.3590 0.7270 3.4090 1.2160 ;
      RECT 2.8630 1.2160 3.4090 1.2660 ;
      RECT 3.8120 0.5270 3.8620 0.6040 ;
      RECT 3.2790 0.4770 3.8620 0.5270 ;
      RECT 2.0060 0.7730 2.7610 0.8230 ;
      RECT 2.5590 0.8230 2.6090 1.1660 ;
      RECT 2.7110 0.8230 2.7610 1.3800 ;
      RECT 2.7110 0.5020 2.7610 0.7730 ;
      RECT 2.5590 0.4520 2.7610 0.5020 ;
      RECT 2.7110 0.3000 2.7610 0.4520 ;
      RECT 2.5590 0.3000 2.6090 0.4520 ;
      RECT 0.8870 1.2020 1.6970 1.2520 ;
      RECT 1.6470 0.7760 1.6970 1.2020 ;
      RECT 1.6470 0.7260 1.7370 0.7760 ;
      RECT 1.6870 0.5760 1.7370 0.7260 ;
      RECT 1.6470 0.5260 1.7370 0.5760 ;
      RECT 1.6470 0.4300 1.6970 0.5260 ;
      RECT 0.8870 1.0970 0.9370 1.2020 ;
      RECT 0.8470 1.0470 0.9370 1.0970 ;
      RECT 0.8470 0.7520 1.0060 0.8020 ;
      RECT 0.9560 0.4930 1.0060 0.7520 ;
      RECT 0.8710 0.4430 1.0060 0.4930 ;
      RECT 0.8470 0.8020 0.8970 1.0470 ;
      RECT 2.1630 0.1540 2.9070 0.2010 ;
      RECT 2.1630 0.1510 3.0050 0.1540 ;
      RECT 2.8570 0.1040 3.0050 0.1510 ;
      RECT 3.5230 0.6770 3.6130 0.7270 ;
      RECT 3.5230 0.7270 3.5730 1.3160 ;
      RECT 2.8110 1.3160 3.5730 1.3660 ;
      RECT 2.8110 1.3660 2.8610 1.5280 ;
      RECT 2.5670 1.5280 2.8610 1.5780 ;
      RECT 2.5670 1.2660 2.6170 1.5280 ;
      RECT 2.4030 1.0440 2.4530 1.2160 ;
      RECT 2.1630 0.9940 2.4530 1.0440 ;
      RECT 2.4030 1.2160 2.6170 1.2660 ;
      RECT 1.7990 0.5730 2.5490 0.6230 ;
      RECT 1.9510 0.4300 2.0010 0.5730 ;
      RECT 1.7990 0.6230 1.8490 1.1960 ;
      RECT 1.7990 0.4300 1.8490 0.5730 ;
      RECT 1.7990 1.1960 2.0010 1.2460 ;
      RECT 1.9510 1.0720 2.0010 1.1960 ;
      RECT 0.4910 1.4490 0.8770 1.4990 ;
      RECT 3.3280 0.1540 3.3780 0.3040 ;
      RECT 2.9750 0.3040 3.3780 0.3540 ;
      RECT 3.2270 0.1040 3.4610 0.1540 ;
      RECT 2.9750 0.3540 3.0250 0.8080 ;
      RECT 2.9750 0.8080 3.0650 0.8580 ;
      RECT 3.0150 0.8580 3.0650 1.1660 ;
      RECT 1.8990 0.6730 2.2450 0.7230 ;
      RECT 1.8990 0.8800 2.1010 0.9300 ;
      RECT 1.8990 0.7230 1.9490 0.8800 ;
      RECT 2.0510 0.9300 2.1010 1.3170 ;
      RECT 1.7590 1.3170 2.1010 1.3670 ;
      RECT 1.7590 1.3670 1.8090 1.5280 ;
      RECT 1.5550 1.5280 1.8090 1.5780 ;
      RECT 1.0990 0.6260 1.4850 0.6760 ;
      RECT 1.1910 0.6760 1.2410 1.1520 ;
      RECT 1.1910 0.4010 1.2410 0.6260 ;
    LAYER PO ;
      RECT 2.1890 0.9660 2.2190 1.6060 ;
      RECT 1.2770 0.0760 1.3070 1.6060 ;
      RECT 2.3410 0.0760 2.3710 1.6060 ;
      RECT 0.8210 0.8700 0.8510 1.6060 ;
      RECT 1.7330 0.0760 1.7630 0.5970 ;
      RECT 2.7970 1.0320 2.8270 1.6060 ;
      RECT 0.5170 0.0760 0.5470 1.6060 ;
      RECT 3.5570 0.0760 3.5870 0.7550 ;
      RECT 3.7090 0.0760 3.7390 1.6060 ;
      RECT 0.8210 0.0760 0.8510 0.6510 ;
      RECT 4.6210 0.0760 4.6510 1.6060 ;
      RECT 1.7330 0.9200 1.7630 1.6060 ;
      RECT 3.8610 0.0760 3.8910 1.6060 ;
      RECT 1.5810 0.0760 1.6110 1.6060 ;
      RECT 4.3170 0.0760 4.3470 1.6060 ;
      RECT 4.1650 0.0760 4.1950 1.6060 ;
      RECT 4.4690 0.0760 4.4990 1.6060 ;
      RECT 4.0130 0.0760 4.0430 1.6060 ;
      RECT 2.0370 0.0760 2.0670 1.6060 ;
      RECT 1.4290 0.0760 1.4590 1.6060 ;
      RECT 2.4930 0.0760 2.5230 1.6060 ;
      RECT 3.5570 1.1320 3.5870 1.6060 ;
      RECT 2.1890 0.0760 2.2190 0.7510 ;
      RECT 3.1010 0.0760 3.1310 1.6060 ;
      RECT 3.4050 0.0760 3.4350 1.6060 ;
      RECT 1.8850 0.0760 1.9150 1.6060 ;
      RECT 3.2530 0.0760 3.2830 1.6060 ;
      RECT 1.1250 0.0760 1.1550 1.6060 ;
      RECT 2.7970 0.0760 2.8270 0.5970 ;
      RECT 2.6450 0.0760 2.6750 1.6060 ;
      RECT 0.6690 0.0760 0.6990 0.5970 ;
      RECT 0.6690 0.8160 0.6990 1.6060 ;
      RECT 2.9490 0.0760 2.9790 1.6060 ;
      RECT 0.9730 0.0760 1.0030 1.6060 ;
      RECT 0.2130 0.0760 0.2430 1.6060 ;
      RECT 0.3650 0.0760 0.3950 1.6060 ;
  END
END DFFSSRX2_LVT

MACRO DFFX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.952 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.9520 0.0300 ;
        RECT 0.5860 0.0300 0.6360 0.1960 ;
        RECT 1.7990 0.0300 1.8490 0.1990 ;
        RECT 0.2790 0.0300 0.3290 0.4190 ;
        RECT 3.4710 0.0300 3.5210 0.2200 ;
        RECT 3.1670 0.0300 3.2170 0.3300 ;
        RECT 0.5860 0.1960 0.9370 0.2460 ;
        RECT 1.7990 0.1990 2.0240 0.2490 ;
        RECT 2.6950 0.3300 3.2330 0.3800 ;
        RECT 0.8870 0.2460 0.9370 0.4500 ;
        RECT 0.7350 0.2460 0.7850 0.4500 ;
        RECT 1.7990 0.2490 1.8490 0.3730 ;
    END
  END VSS

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.7450 1.1610 3.8560 1.2210 ;
        RECT 3.6230 1.2210 3.8560 1.2710 ;
        RECT 3.8050 0.2040 3.8550 1.1610 ;
        RECT 3.6230 1.2710 3.6730 1.5460 ;
        RECT 3.6070 0.1540 3.8550 0.2040 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.9520 1.7020 ;
        RECT 0.2790 1.0330 0.3290 1.6420 ;
        RECT 3.4710 0.9470 3.5210 1.6420 ;
        RECT 0.8870 1.3540 0.9370 1.6420 ;
        RECT 2.6390 1.3580 2.6890 1.6420 ;
        RECT 1.9750 1.3280 2.0250 1.6420 ;
        RECT 3.2070 1.3580 3.2570 1.6420 ;
        RECT 0.7350 1.3040 0.9370 1.3540 ;
        RECT 2.6390 1.3080 2.7770 1.3580 ;
        RECT 1.7820 1.2780 2.0250 1.3280 ;
        RECT 3.1490 1.3080 3.2570 1.3580 ;
        RECT 0.7350 1.0880 0.7850 1.3040 ;
        RECT 0.8870 1.1010 0.9370 1.3040 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.3590 0.6800 ;
        RECT 0.2490 0.6800 0.4210 0.7300 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.4240 0.7250 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.5930 1.0090 3.7030 1.1190 ;
        RECT 3.6530 0.8540 3.7030 1.0090 ;
        RECT 3.3190 0.8040 3.7030 0.8540 ;
        RECT 3.3190 0.8540 3.3690 1.5460 ;
        RECT 3.6530 0.3590 3.7030 0.8040 ;
        RECT 3.3190 0.3090 3.7030 0.3590 ;
        RECT 3.3190 0.1480 3.3690 0.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 4.0670 1.7730 ;
    LAYER M1 ;
      RECT 1.1910 0.2990 1.2810 0.3810 ;
      RECT 1.2150 0.3810 1.2650 0.9880 ;
      RECT 1.1910 1.0380 1.2410 1.3140 ;
      RECT 0.4310 0.9880 1.2650 1.0380 ;
      RECT 0.4310 1.0380 0.4810 1.2160 ;
      RECT 0.4310 0.8290 0.4810 0.9880 ;
      RECT 0.4310 0.5790 0.5210 0.6290 ;
      RECT 0.4310 0.4550 0.4810 0.5790 ;
      RECT 0.4310 0.7800 0.5210 0.8290 ;
      RECT 0.4710 0.6290 0.5210 0.7800 ;
      RECT 2.7870 0.0880 2.8370 0.2300 ;
      RECT 2.1150 0.2300 2.8370 0.2800 ;
      RECT 2.3150 0.1780 2.3970 0.2300 ;
      RECT 2.1150 0.2800 2.1650 0.3140 ;
      RECT 1.9640 0.3140 2.1650 0.3640 ;
      RECT 1.9640 0.3640 2.0140 0.5400 ;
      RECT 1.7070 0.5400 2.0140 0.5900 ;
      RECT 1.3430 0.6400 2.0930 0.6900 ;
      RECT 1.3430 0.6900 1.3930 1.1580 ;
      RECT 1.3430 0.4840 1.3930 0.6400 ;
      RECT 1.3430 1.1580 1.5610 1.2080 ;
      RECT 1.3430 0.4340 1.5610 0.4840 ;
      RECT 1.3430 1.2080 1.3930 1.3140 ;
      RECT 1.3430 0.3550 1.3930 0.4340 ;
      RECT 3.5470 0.4880 3.5970 0.7040 ;
      RECT 2.4070 0.4380 3.5970 0.4880 ;
      RECT 3.2070 0.7040 3.5970 0.7540 ;
      RECT 3.2070 0.7540 3.2570 1.2080 ;
      RECT 2.8470 1.2080 3.2570 1.2580 ;
      RECT 2.4070 0.4880 2.4570 1.1650 ;
      RECT 2.7100 0.4880 2.7600 0.6990 ;
      RECT 2.6190 0.6990 2.7600 0.7490 ;
      RECT 1.7070 0.7580 2.2290 0.8080 ;
      RECT 2.1790 0.5870 2.2290 0.7580 ;
      RECT 1.5500 1.0010 2.3450 1.0510 ;
      RECT 2.2950 0.4700 2.3450 1.0010 ;
      RECT 2.2550 1.0510 2.3050 1.3080 ;
      RECT 2.0720 0.4200 2.3450 0.4700 ;
      RECT 2.1030 1.3080 2.3050 1.3580 ;
      RECT 2.2550 0.3710 2.3050 0.4200 ;
      RECT 2.1030 1.1660 2.1530 1.3080 ;
      RECT 2.8240 0.6040 3.4610 0.6540 ;
      RECT 2.8240 0.6540 2.8740 0.9780 ;
      RECT 2.5190 0.9780 2.8740 1.0270 ;
      RECT 2.5420 1.0270 2.8740 1.0280 ;
      RECT 2.5190 0.5880 2.5690 0.9780 ;
      RECT 2.8240 1.0280 2.8740 1.0290 ;
      RECT 2.5190 0.5380 2.6490 0.5880 ;
      RECT 2.7700 1.5210 3.1570 1.5710 ;
      RECT 1.4190 1.4780 1.7890 1.5280 ;
      RECT 1.4190 1.5280 1.4690 1.5650 ;
      RECT 1.0990 1.5260 1.3170 1.5760 ;
      RECT 1.2670 1.4280 1.3170 1.5260 ;
      RECT 1.2670 1.3780 1.9250 1.4280 ;
      RECT 1.8750 1.4280 1.9250 1.5840 ;
      RECT 0.5830 0.6180 1.0290 0.6680 ;
      RECT 0.5830 0.6680 0.6330 0.9140 ;
      RECT 0.5830 0.4220 0.6330 0.6180 ;
      RECT 1.0390 0.5180 1.1650 0.5680 ;
      RECT 1.0390 0.3940 1.0890 0.5180 ;
      RECT 1.1150 0.5680 1.1650 0.7180 ;
      RECT 1.0390 0.7180 1.1650 0.7680 ;
      RECT 1.0390 0.7680 1.0890 0.9140 ;
      RECT 2.9340 0.7090 3.1570 0.7590 ;
      RECT 2.5310 1.1490 2.5810 1.2720 ;
      RECT 2.3550 1.2720 2.5810 1.3220 ;
      RECT 2.3550 1.3220 2.4050 1.5220 ;
      RECT 2.1630 1.5220 2.4050 1.5720 ;
      RECT 2.9340 0.7590 2.9840 1.0990 ;
      RECT 2.5310 1.0990 2.9840 1.1490 ;
      RECT 0.7950 0.0960 1.4910 0.1460 ;
    LAYER PO ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 1.2770 0.0680 1.3070 0.5420 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 1.2770 0.9900 1.3070 1.6060 ;
      RECT 3.1010 0.0680 3.1310 0.7870 ;
      RECT 1.7330 0.0680 1.7630 0.6180 ;
      RECT 2.3410 0.8820 2.3710 1.6060 ;
      RECT 3.1010 1.0120 3.1310 1.6060 ;
      RECT 2.3410 0.0680 2.3710 0.6220 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 1.7330 0.7300 1.7630 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 3.7090 0.0680 3.7390 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
  END
END DFFX1_LVT

MACRO DFFX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.256 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0490 0.0970 4.1590 0.2070 ;
        RECT 4.0910 0.2070 4.1410 0.2700 ;
        RECT 3.7750 0.2700 4.1410 0.3200 ;
        RECT 3.7750 0.1480 3.8250 0.2700 ;
        RECT 4.0910 0.3200 4.1410 0.9180 ;
        RECT 3.7750 0.9180 4.1410 0.9680 ;
        RECT 3.7750 0.9680 3.8250 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4710 0.1480 3.5210 0.3940 ;
        RECT 3.4710 0.3940 4.0170 0.4440 ;
        RECT 3.8970 0.4440 4.0170 0.5110 ;
        RECT 3.9670 0.5110 4.0170 0.8040 ;
        RECT 3.4710 0.8040 4.0170 0.8540 ;
        RECT 3.4710 0.8540 3.5210 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.2560 0.0300 ;
        RECT 0.5860 0.0300 0.6360 0.1960 ;
        RECT 1.7990 0.0300 1.8490 0.1990 ;
        RECT 3.3190 0.0300 3.3690 0.4080 ;
        RECT 3.9270 0.0300 3.9770 0.2200 ;
        RECT 0.2790 0.0300 0.3290 0.4190 ;
        RECT 3.6230 0.0300 3.6730 0.3190 ;
        RECT 3.1670 0.0300 3.2170 0.3300 ;
        RECT 0.5860 0.1960 0.9370 0.2460 ;
        RECT 1.7990 0.1990 2.0240 0.2490 ;
        RECT 2.6950 0.3300 3.2330 0.3800 ;
        RECT 0.8870 0.2460 0.9370 0.4500 ;
        RECT 0.7350 0.2460 0.7850 0.4500 ;
        RECT 1.7990 0.2490 1.8490 0.3730 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.2560 1.7020 ;
        RECT 0.2790 1.0330 0.3290 1.6420 ;
        RECT 3.3190 0.9120 3.3690 1.6420 ;
        RECT 3.9270 1.0520 3.9770 1.6420 ;
        RECT 3.6230 0.9600 3.6730 1.6420 ;
        RECT 0.8870 1.3540 0.9370 1.6420 ;
        RECT 1.9750 1.3280 2.0250 1.6420 ;
        RECT 3.2070 1.3580 3.2570 1.6420 ;
        RECT 2.6390 1.3580 2.6890 1.6420 ;
        RECT 0.7350 1.3040 0.9370 1.3540 ;
        RECT 1.7820 1.2780 2.0250 1.3280 ;
        RECT 3.1490 1.3080 3.2570 1.3580 ;
        RECT 2.6390 1.3080 2.7770 1.3580 ;
        RECT 0.7350 1.0880 0.7850 1.3040 ;
        RECT 0.8870 1.1010 0.9370 1.3040 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.3590 0.6800 ;
        RECT 0.2490 0.6800 0.4210 0.7300 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.4240 0.7250 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 4.3710 1.7730 ;
    LAYER M1 ;
      RECT 1.1910 0.2990 1.2810 0.3810 ;
      RECT 1.2150 0.3810 1.2650 0.9880 ;
      RECT 1.1910 1.0380 1.2410 1.3140 ;
      RECT 0.4310 0.9880 1.2650 1.0380 ;
      RECT 0.4310 1.0380 0.4810 1.2160 ;
      RECT 0.4310 0.8290 0.4810 0.9880 ;
      RECT 0.4310 0.5790 0.5210 0.6290 ;
      RECT 0.4310 0.4550 0.4810 0.5790 ;
      RECT 0.4310 0.7800 0.5210 0.8290 ;
      RECT 0.4710 0.6290 0.5210 0.7800 ;
      RECT 2.7870 0.0880 2.8370 0.2300 ;
      RECT 2.1150 0.2300 2.8370 0.2800 ;
      RECT 2.3150 0.1780 2.3970 0.2300 ;
      RECT 2.1150 0.2800 2.1650 0.3140 ;
      RECT 1.9640 0.3140 2.1650 0.3640 ;
      RECT 1.9640 0.3640 2.0140 0.5400 ;
      RECT 1.7070 0.5400 2.0140 0.5900 ;
      RECT 1.3430 0.6400 2.0930 0.6900 ;
      RECT 1.3430 0.6900 1.3930 1.1580 ;
      RECT 1.3430 0.4840 1.3930 0.6400 ;
      RECT 1.3430 1.1580 1.5610 1.2080 ;
      RECT 1.3430 0.4340 1.5610 0.4840 ;
      RECT 1.3430 1.2080 1.3930 1.3140 ;
      RECT 1.3430 0.3550 1.3930 0.4340 ;
      RECT 3.6800 0.6040 3.9170 0.6540 ;
      RECT 2.7100 0.5440 2.7600 0.6990 ;
      RECT 2.7100 0.4880 2.7600 0.4940 ;
      RECT 3.2070 0.7540 3.2570 1.2080 ;
      RECT 2.6190 0.6990 2.7600 0.7490 ;
      RECT 2.4070 0.4380 2.7600 0.4880 ;
      RECT 2.8470 1.2080 3.2570 1.2580 ;
      RECT 2.4070 0.4880 2.4570 1.1650 ;
      RECT 3.6800 0.5440 3.7300 0.6040 ;
      RECT 3.6800 0.6540 3.7300 0.7040 ;
      RECT 3.2070 0.7040 3.7300 0.7540 ;
      RECT 2.7100 0.4940 3.7300 0.5440 ;
      RECT 1.7070 0.7580 2.2290 0.8080 ;
      RECT 2.1790 0.5870 2.2290 0.7580 ;
      RECT 1.5500 1.0010 2.3450 1.0510 ;
      RECT 2.2950 0.4700 2.3450 1.0010 ;
      RECT 2.2550 1.0510 2.3050 1.3080 ;
      RECT 2.0720 0.4200 2.3450 0.4700 ;
      RECT 2.1030 1.3080 2.3050 1.3580 ;
      RECT 2.2550 0.3710 2.3050 0.4200 ;
      RECT 2.1030 1.1660 2.1530 1.3080 ;
      RECT 2.7700 1.5210 3.1570 1.5710 ;
      RECT 1.4190 1.4780 1.7890 1.5280 ;
      RECT 1.4190 1.5280 1.4690 1.5650 ;
      RECT 1.0990 1.5260 1.3170 1.5760 ;
      RECT 1.2670 1.4280 1.3170 1.5260 ;
      RECT 1.2670 1.3780 1.9250 1.4280 ;
      RECT 1.8750 1.4280 1.9250 1.5840 ;
      RECT 0.5830 0.6180 1.0290 0.6680 ;
      RECT 0.5830 0.6680 0.6330 0.9140 ;
      RECT 0.5830 0.4220 0.6330 0.6180 ;
      RECT 1.0390 0.5180 1.1650 0.5680 ;
      RECT 1.0390 0.3940 1.0890 0.5180 ;
      RECT 1.1150 0.5680 1.1650 0.7180 ;
      RECT 1.0390 0.7180 1.1650 0.7680 ;
      RECT 1.0390 0.7680 1.0890 0.9140 ;
      RECT 2.8240 0.6040 3.6130 0.6540 ;
      RECT 2.8240 0.6540 2.8740 0.9780 ;
      RECT 2.5190 0.9780 2.8740 1.0270 ;
      RECT 2.5190 0.5880 2.5690 0.9780 ;
      RECT 2.5420 1.0270 2.8740 1.0280 ;
      RECT 2.5190 0.5380 2.6250 0.5880 ;
      RECT 2.8240 1.0280 2.8740 1.0290 ;
      RECT 2.9340 0.7090 3.1570 0.7590 ;
      RECT 2.5310 1.1490 2.5810 1.2720 ;
      RECT 2.3550 1.2720 2.5810 1.3220 ;
      RECT 2.3550 1.3220 2.4050 1.5220 ;
      RECT 2.1630 1.5220 2.4050 1.5720 ;
      RECT 2.9340 0.7590 2.9840 1.0990 ;
      RECT 2.5310 1.0990 2.9840 1.1490 ;
      RECT 0.7950 0.0960 1.4910 0.1460 ;
    LAYER PO ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 3.7090 0.0680 3.7390 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 1.2770 0.0680 1.3070 0.5420 ;
      RECT 1.2770 0.9900 1.3070 1.6060 ;
      RECT 3.1010 0.0680 3.1310 0.7870 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 1.7330 0.0680 1.7630 0.6180 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 2.3410 0.8820 2.3710 1.6060 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 3.1010 1.0120 3.1310 1.6060 ;
      RECT 2.3410 0.0680 2.3710 0.6220 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 1.7330 0.7300 1.7630 1.6060 ;
  END
END DFFX2_LVT

MACRO DHFILLH2_LVT
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.304 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 0.3040 0.0300 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 0.3040 3.3740 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 0.3040 1.7020 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1150 2.3510 0.4190 3.4450 ;
      RECT -0.1150 -0.1010 0.4190 0.9930 ;
    LAYER PO ;
      RECT 0.0610 1.7900 0.0910 3.2680 ;
      RECT 0.2130 1.7890 0.2430 3.2670 ;
      RECT 0.2130 0.1170 0.2430 1.5960 ;
      RECT 0.0610 0.1180 0.0910 1.5960 ;
  END
END DHFILLH2_LVT

MACRO DHFILLHL2_LVT
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.304 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 0.3040 1.7020 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 0.3040 0.0300 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 0.3040 3.3740 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 0.4190 2.6650 ;
    LAYER PO ;
      RECT 0.0610 0.1190 0.0910 1.5970 ;
      RECT 0.2130 0.1180 0.2430 1.5970 ;
      RECT 0.0610 1.7910 0.0910 3.2690 ;
      RECT 0.2130 1.7900 0.2430 3.2680 ;
  END
END DHFILLHL2_LVT

MACRO DHFILLHLHLS11_LVT
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.672 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.6720 0.0300 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 1.6720 3.3740 ;
    END
  END VDDH

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.6720 1.7020 ;
    END
  END VSS

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 3.0100 1.6720 3.0700 ;
        RECT 0.8080 2.5310 0.8640 3.0100 ;
    END
  END VDDL
  OBS
    LAYER NWELL ;
      RECT -0.1150 -0.1010 1.7870 0.9930 ;
      RECT -0.1150 2.3510 1.7870 3.4450 ;
    LAYER PO ;
      RECT 1.4290 0.1070 1.4590 1.5850 ;
      RECT 1.5810 0.1060 1.6110 1.5850 ;
      RECT 1.5810 1.7780 1.6110 3.2560 ;
      RECT 1.4290 1.7790 1.4590 3.2570 ;
      RECT 1.2770 1.7780 1.3070 3.2560 ;
      RECT 1.2770 0.1060 1.3070 1.5850 ;
      RECT 1.1250 0.1070 1.1550 1.5850 ;
      RECT 1.1250 1.7790 1.1550 3.2570 ;
      RECT 0.3650 1.7790 0.3950 3.2570 ;
      RECT 0.5170 1.7780 0.5470 3.2560 ;
      RECT 0.5170 0.1060 0.5470 1.5850 ;
      RECT 0.0610 1.7810 0.0910 3.2590 ;
      RECT 0.0610 0.1090 0.0910 1.5870 ;
      RECT 0.3650 0.1070 0.3950 1.5850 ;
      RECT 0.2130 0.1080 0.2430 1.5870 ;
      RECT 0.2130 1.7800 0.2430 3.2580 ;
  END
END DHFILLHLHLS11_LVT

MACRO FADDX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.888 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6430 0.5940 1.8100 0.6440 ;
        RECT 0.7050 0.6440 0.8150 0.6630 ;
        RECT 0.7050 0.5530 0.8150 0.5940 ;
    END
    ANTENNAGATEAREA 0.081 ;
  END CI

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8610 1.1610 0.9920 1.2710 ;
        RECT 0.8610 0.8760 0.9110 1.1610 ;
        RECT 0.3390 0.8260 2.0770 0.8760 ;
        RECT 2.0270 0.8760 2.0770 0.8920 ;
        RECT 2.0270 0.8100 2.0770 0.8260 ;
    END
    ANTENNAGATEAREA 0.108 ;
  END A

  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5590 0.8420 2.6330 0.8570 ;
        RECT 2.5830 0.5610 2.6330 0.8420 ;
        RECT 2.5590 0.8570 2.7910 0.9670 ;
        RECT 2.5590 0.4790 2.6330 0.5610 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END CO

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 0.5530 0.5110 0.7130 ;
        RECT 0.4010 0.7130 1.9490 0.7630 ;
    END
    ANTENNAGATEAREA 0.108 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.0040 1.6420 2.8880 1.7020 ;
        RECT 2.1030 1.4400 2.1530 1.6420 ;
        RECT 1.3430 1.4340 1.3930 1.6420 ;
        RECT 1.0390 1.4380 1.0890 1.6420 ;
        RECT 0.4310 1.4380 0.4810 1.6420 ;
        RECT 2.4070 1.3230 2.4570 1.6420 ;
    END
  END VDD

  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2310 0.5610 2.2810 1.0090 ;
        RECT 2.2310 1.0090 2.4870 1.1190 ;
        RECT 2.2310 0.4790 2.3050 0.5610 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END S

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.8880 0.0300 ;
        RECT 0.4310 0.0300 0.4810 0.2030 ;
        RECT 2.1030 0.0300 2.1530 0.2030 ;
        RECT 2.4070 0.0300 2.4570 0.2030 ;
        RECT 1.0390 0.0300 1.0890 0.2370 ;
        RECT 1.0390 0.2370 1.4090 0.2870 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 3.0030 1.7730 ;
    LAYER M1 ;
      RECT 2.4550 0.6240 2.5330 0.7140 ;
      RECT 1.5310 0.2530 2.5050 0.3030 ;
      RECT 2.4550 0.3030 2.5050 0.6240 ;
      RECT 2.4550 0.7140 2.5050 0.7290 ;
      RECT 1.5310 0.3030 1.5810 0.3550 ;
      RECT 0.2390 0.3550 1.5810 0.4050 ;
      RECT 1.5310 0.4050 1.5810 0.4750 ;
      RECT 1.5310 0.4750 1.6370 0.5250 ;
      RECT 0.2390 1.0570 0.8010 1.1070 ;
      RECT 0.2390 0.4050 0.2890 1.0570 ;
      RECT 1.6310 0.3550 2.4050 0.4050 ;
      RECT 2.3550 0.7140 2.4050 0.7290 ;
      RECT 1.6310 1.0790 2.1810 1.1290 ;
      RECT 2.3310 0.6240 2.4050 0.7140 ;
      RECT 2.3550 0.4050 2.4050 0.6240 ;
      RECT 2.1310 0.4050 2.1810 1.0790 ;
      RECT 1.1750 0.1370 1.5610 0.1870 ;
      RECT 0.2630 1.2230 0.6490 1.2730 ;
      RECT 0.2630 0.2550 0.6490 0.3050 ;
      RECT 1.1750 1.2230 1.5610 1.2730 ;
    LAYER PO ;
      RECT 2.1890 0.0710 2.2190 1.6090 ;
      RECT 0.5170 0.0710 0.5470 1.6090 ;
      RECT 0.6690 0.0710 0.6990 1.6090 ;
      RECT 1.1250 0.0710 1.1550 1.6090 ;
      RECT 1.7330 0.0710 1.7630 1.6090 ;
      RECT 2.6450 0.0710 2.6750 1.6090 ;
      RECT 2.7970 0.0710 2.8270 1.6090 ;
      RECT 1.4290 0.0710 1.4590 1.6090 ;
      RECT 0.2130 0.0710 0.2430 1.6090 ;
      RECT 1.2770 0.0710 1.3070 1.6090 ;
      RECT 0.9730 0.0670 1.0030 1.6090 ;
      RECT 0.0610 0.0710 0.0910 1.6090 ;
      RECT 1.5810 0.0710 1.6110 1.6090 ;
      RECT 2.4930 0.0710 2.5230 1.6090 ;
      RECT 2.3410 0.0710 2.3710 1.6090 ;
      RECT 0.3650 0.0710 0.3950 1.6090 ;
      RECT 0.8210 0.0710 0.8510 1.6090 ;
      RECT 2.0370 0.0710 2.0670 1.6090 ;
      RECT 1.8850 0.0710 1.9150 1.6090 ;
  END
END FADDX1_LVT

MACRO FADDX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.192 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6430 0.5470 1.8100 0.5970 ;
        RECT 0.6700 0.5970 0.8430 0.6650 ;
    END
    ANTENNAGATEAREA 0.081 ;
  END CI

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8010 1.1610 0.9670 1.2710 ;
        RECT 0.8610 0.8730 0.9110 1.1610 ;
        RECT 0.3390 0.8230 2.0770 0.8730 ;
        RECT 2.0270 0.8730 2.0770 0.8890 ;
        RECT 2.0270 0.8070 2.0770 0.8230 ;
    END
    ANTENNAGATEAREA 0.108 ;
  END A

  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.7110 0.4950 2.9370 0.5450 ;
        RECT 2.7110 0.4790 2.7610 0.4950 ;
        RECT 2.7110 0.5450 2.7610 0.5610 ;
        RECT 2.8870 0.5450 2.9370 0.8420 ;
        RECT 2.8870 0.4790 2.9370 0.4950 ;
        RECT 2.7110 0.8420 2.9420 0.8570 ;
        RECT 2.7110 0.8570 3.0950 0.8920 ;
        RECT 2.7110 0.8920 2.7610 0.9290 ;
        RECT 2.8870 0.8920 3.0950 0.9670 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END CO

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 0.5530 0.5110 0.6650 ;
        RECT 0.4280 0.6650 0.4840 0.7230 ;
        RECT 0.3450 0.7230 1.9490 0.7730 ;
    END
    ANTENNAGATEAREA 0.108 ;
  END B

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.1920 1.7020 ;
        RECT 2.1030 1.3230 2.1530 1.6420 ;
        RECT 1.3430 1.3230 1.3930 1.6420 ;
        RECT 1.0390 1.3230 1.0890 1.6420 ;
        RECT 0.4310 1.3230 0.4810 1.6420 ;
        RECT 2.8630 1.3230 2.9130 1.6420 ;
        RECT 2.2550 1.3230 2.3050 1.6420 ;
        RECT 2.5590 1.3230 2.6090 1.6420 ;
    END
  END VDD

  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2310 0.4790 2.4570 0.5290 ;
        RECT 2.2310 0.5290 2.2810 1.0090 ;
        RECT 2.4070 0.5290 2.4570 0.5610 ;
        RECT 2.2310 1.0090 2.4870 1.1190 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END S

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.1920 0.0300 ;
        RECT 0.3710 0.0300 0.4210 0.1370 ;
        RECT 2.5590 0.0300 2.6090 0.1470 ;
        RECT 1.0390 0.0300 1.0890 0.2370 ;
        RECT 0.3710 0.1370 0.5160 0.1870 ;
        RECT 2.0850 0.1470 2.9340 0.1970 ;
        RECT 1.0390 0.2370 1.4090 0.2870 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 3.3070 1.7730 ;
    LAYER M1 ;
      RECT 2.6070 0.6210 2.8370 0.7110 ;
      RECT 2.6070 0.7110 2.6570 0.7290 ;
      RECT 2.6070 0.2970 2.6570 0.6210 ;
      RECT 1.5310 0.2470 2.6570 0.2970 ;
      RECT 1.5310 0.2970 1.5810 0.3550 ;
      RECT 0.2390 0.3550 1.5810 0.4050 ;
      RECT 1.5310 0.4050 1.5810 0.4470 ;
      RECT 1.5310 0.4470 1.6370 0.4970 ;
      RECT 0.2390 1.0570 0.8010 1.1070 ;
      RECT 0.2390 0.4050 0.2890 1.0570 ;
      RECT 2.5070 0.7110 2.5570 0.7290 ;
      RECT 1.6310 0.3470 2.5570 0.3970 ;
      RECT 2.3310 0.6210 2.5570 0.7110 ;
      RECT 2.5070 0.3970 2.5570 0.6210 ;
      RECT 1.6310 1.0790 2.1810 1.1290 ;
      RECT 2.1310 0.3970 2.1810 1.0790 ;
      RECT 1.1750 0.1370 1.5610 0.1870 ;
      RECT 0.2630 1.2230 0.6490 1.2730 ;
      RECT 0.2630 0.2370 0.6490 0.2870 ;
      RECT 1.1750 1.2230 1.5610 1.2730 ;
    LAYER PO ;
      RECT 2.1890 0.0710 2.2190 1.6090 ;
      RECT 0.5170 0.0710 0.5470 1.6090 ;
      RECT 0.6690 0.0710 0.6990 1.6090 ;
      RECT 1.1250 0.0710 1.1550 1.6090 ;
      RECT 1.7330 0.0710 1.7630 1.6090 ;
      RECT 2.6450 0.0710 2.6750 1.6090 ;
      RECT 2.7970 0.0710 2.8270 1.6090 ;
      RECT 1.4290 0.0710 1.4590 1.6090 ;
      RECT 0.2130 0.0710 0.2430 1.6090 ;
      RECT 1.2770 0.0710 1.3070 1.6090 ;
      RECT 0.9730 0.0670 1.0030 1.6090 ;
      RECT 0.0610 0.0710 0.0910 1.6090 ;
      RECT 1.5810 0.0710 1.6110 1.6090 ;
      RECT 2.4930 0.0710 2.5230 1.6090 ;
      RECT 2.3410 0.0710 2.3710 1.6090 ;
      RECT 3.1010 0.0710 3.1310 1.6090 ;
      RECT 0.3650 0.0710 0.3950 1.6090 ;
      RECT 0.8210 0.0710 0.8510 1.6090 ;
      RECT 2.9490 0.0710 2.9790 1.6090 ;
      RECT 2.0370 0.0710 2.0670 1.6090 ;
      RECT 1.8850 0.0710 1.9150 1.6090 ;
  END
END FADDX2_LVT

MACRO FOOT2X16_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.6 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VSSG
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.7500 1.1750 0.9940 1.2570 ;
        RECT 0.8860 1.2570 0.9360 1.5340 ;
        RECT 0.8710 1.5340 6.7290 1.5900 ;
    END
  END VSSG

  PIN VSS
    DIRECTION OUTPUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 7.6000 1.7020 ;
        RECT 5.5990 1.7020 5.6490 1.8320 ;
        RECT 6.5110 1.7020 6.5610 1.8320 ;
        RECT 4.9910 1.7020 5.0410 1.8320 ;
        RECT 4.0790 1.7020 4.1290 1.8320 ;
        RECT 2.5590 1.7020 2.6090 1.8320 ;
        RECT 3.4710 1.7020 3.5210 1.8320 ;
        RECT 1.9510 1.7020 2.0010 1.8320 ;
        RECT 1.0390 1.7020 1.0890 1.8320 ;
    END
  END VSS

  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8000 2.1560 0.9670 2.1810 ;
        RECT 0.8000 2.1060 6.8270 2.1560 ;
        RECT 0.8000 2.0710 0.9670 2.1060 ;
    END
    ANTENNAGATEAREA 0.1248 ;
  END SLEEP

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 7.6000 0.0300 ;
        RECT 5.7510 0.0300 5.8010 0.9240 ;
        RECT 6.0550 0.0300 6.1050 0.9240 ;
        RECT 6.3590 0.0300 6.4090 0.9240 ;
        RECT 4.8390 0.0300 4.8890 0.9240 ;
        RECT 4.5350 0.0300 4.5850 0.9240 ;
        RECT 4.2310 0.0300 4.2810 0.9240 ;
        RECT 2.7110 0.0300 2.7610 0.9240 ;
        RECT 3.0150 0.0300 3.0650 0.9240 ;
        RECT 3.3190 0.0300 3.3690 0.9240 ;
        RECT 1.7990 0.0300 1.8490 0.9240 ;
        RECT 1.4950 0.0300 1.5450 0.9240 ;
        RECT 1.1910 0.0300 1.2410 0.9240 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 7.6000 3.3740 ;
        RECT 0.8870 2.4720 0.9370 3.3140 ;
    END
  END VDD

  PIN SLEEPOUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.1770 1.2000 6.2870 1.2710 ;
        RECT 6.2070 1.2710 6.2570 1.4840 ;
        RECT 1.3430 1.1610 6.2870 1.2000 ;
        RECT 1.3430 1.2000 1.3930 1.4840 ;
        RECT 2.8630 1.2000 2.9130 1.4840 ;
        RECT 1.6470 1.2000 1.6970 1.4840 ;
        RECT 4.3830 1.2000 4.4330 1.4840 ;
        RECT 3.1670 1.2000 3.2170 1.4840 ;
        RECT 4.6870 1.2000 4.7370 1.4840 ;
        RECT 1.3430 1.1500 6.2570 1.1610 ;
        RECT 5.9030 1.2000 5.9530 1.4840 ;
        RECT 1.3430 0.1980 1.3930 1.1500 ;
        RECT 2.8630 0.1980 2.9130 1.1500 ;
        RECT 1.6470 0.1980 1.6970 1.1500 ;
        RECT 4.3830 0.1980 4.4330 1.1500 ;
        RECT 3.1670 0.1980 3.2170 1.1500 ;
        RECT 4.6870 0.1980 4.7370 1.1500 ;
        RECT 5.9030 0.1980 5.9530 1.1500 ;
        RECT 6.2070 0.1980 6.2570 1.1500 ;
    END
    ANTENNADIFFAREA 1.1904 ;
  END SLEEPOUT
  OBS
    LAYER PO ;
      RECT 2.6450 0.0510 2.6750 0.9710 ;
      RECT 3.4050 0.0510 3.4350 0.9710 ;
      RECT 2.3410 1.3510 2.3710 2.1670 ;
      RECT 2.6450 1.3510 2.6750 1.9790 ;
      RECT 2.4930 1.3510 2.5230 1.9790 ;
      RECT 3.4050 1.3510 3.4350 1.9790 ;
      RECT 3.5570 1.3510 3.5870 1.9790 ;
      RECT 6.7490 1.3510 6.7790 2.1670 ;
      RECT 1.5810 0.0510 1.6110 1.9790 ;
      RECT 1.7330 0.0510 1.7630 1.9790 ;
      RECT 1.8850 0.0510 1.9150 0.9710 ;
      RECT 1.8850 1.3510 1.9150 1.9790 ;
      RECT 2.0370 1.3510 2.0670 1.9790 ;
      RECT 3.7090 1.3510 3.7390 2.1670 ;
      RECT 2.1890 1.3510 2.2190 2.1670 ;
      RECT 0.9730 2.3730 1.0030 3.2930 ;
      RECT 1.4290 0.0510 1.4590 1.9790 ;
      RECT 1.1250 0.0510 1.1550 0.9710 ;
      RECT 0.6690 2.3730 0.6990 3.2930 ;
      RECT 1.2770 0.0510 1.3070 1.9790 ;
      RECT 0.6690 1.3510 0.6990 1.8920 ;
      RECT 0.8210 1.3510 0.8510 3.2930 ;
      RECT 1.1250 1.3510 1.1550 1.9790 ;
      RECT 0.9730 1.3510 1.0030 1.9790 ;
      RECT 2.9490 2.3730 2.9790 3.2930 ;
      RECT 2.1890 2.3730 2.2190 3.2930 ;
      RECT 4.0130 2.3730 4.0430 3.2930 ;
      RECT 4.1650 2.3730 4.1950 3.2930 ;
      RECT 4.3170 2.3730 4.3470 3.2930 ;
      RECT 3.8610 2.3730 3.8910 3.2930 ;
      RECT 3.7090 2.3730 3.7390 3.2930 ;
      RECT 3.5570 2.3730 3.5870 3.2930 ;
      RECT 3.4050 2.3730 3.4350 3.2930 ;
      RECT 3.2530 2.3730 3.2830 3.2930 ;
      RECT 5.5330 2.3730 5.5630 3.2930 ;
      RECT 5.6850 2.3730 5.7150 3.2930 ;
      RECT 5.8370 2.3730 5.8670 3.2930 ;
      RECT 5.9890 2.3730 6.0190 3.2930 ;
      RECT 6.4440 2.3730 6.4750 3.2930 ;
      RECT 6.2930 2.3730 6.3230 3.2930 ;
      RECT 6.1410 2.3730 6.1710 3.2930 ;
      RECT 5.3810 2.3730 5.4110 3.2930 ;
      RECT 7.2050 2.3730 7.2350 3.2930 ;
      RECT 7.3570 2.3730 7.3870 3.2930 ;
      RECT 7.5090 2.3730 7.5390 3.2930 ;
      RECT 7.0530 2.3730 7.0830 3.2930 ;
      RECT 6.9010 2.3730 6.9310 3.2930 ;
      RECT 6.7490 2.3730 6.7790 3.2930 ;
      RECT 6.5970 2.3730 6.6270 3.2930 ;
      RECT 1.7330 2.3730 1.7630 3.2930 ;
      RECT 1.8850 2.3730 1.9150 3.2930 ;
      RECT 2.0370 2.3730 2.0670 3.2930 ;
      RECT 1.5810 2.3730 1.6110 3.2930 ;
      RECT 0.5170 2.3730 0.5470 3.2930 ;
      RECT 0.3650 2.3730 0.3950 3.2930 ;
      RECT 0.2130 2.3730 0.2430 3.2930 ;
      RECT 0.0610 2.3730 0.0910 3.2930 ;
      RECT 1.4290 2.3730 1.4590 3.2930 ;
      RECT 1.2770 2.3730 1.3070 3.2930 ;
      RECT 1.1250 2.3730 1.1550 3.2930 ;
      RECT 7.3570 1.3510 7.3870 1.8920 ;
      RECT 7.2050 1.3510 7.2350 1.8920 ;
      RECT 7.5090 1.3510 7.5390 1.8920 ;
      RECT 7.0530 1.3510 7.0830 1.8920 ;
      RECT 0.5170 1.3510 0.5470 1.8920 ;
      RECT 0.3650 1.3510 0.3950 1.8920 ;
      RECT 0.2130 1.3510 0.2430 1.8920 ;
      RECT 0.0610 1.3510 0.0910 1.8920 ;
      RECT 0.6690 0.0510 0.6990 0.9710 ;
      RECT 0.8210 0.0510 0.8510 0.9710 ;
      RECT 0.9730 0.0510 1.0030 0.9710 ;
      RECT 0.3650 0.0510 0.3950 0.9710 ;
      RECT 0.5170 0.0510 0.5470 0.9710 ;
      RECT 0.2130 0.0510 0.2430 0.9710 ;
      RECT 0.0610 0.0510 0.0910 0.9710 ;
      RECT 2.3410 0.0510 2.3710 0.9710 ;
      RECT 2.4930 0.0510 2.5230 0.9710 ;
      RECT 2.1890 0.0510 2.2190 0.9710 ;
      RECT 2.0370 0.0510 2.0670 0.9710 ;
      RECT 3.5570 0.0510 3.5870 0.9710 ;
      RECT 3.7090 0.0510 3.7390 0.9710 ;
      RECT 4.0130 0.0510 4.0430 0.9710 ;
      RECT 3.8610 0.0510 3.8910 0.9710 ;
      RECT 5.0770 0.0510 5.1070 0.9710 ;
      RECT 5.2290 0.0510 5.2590 0.9710 ;
      RECT 5.5330 0.0510 5.5630 0.9710 ;
      RECT 5.3810 0.0510 5.4110 0.9710 ;
      RECT 6.5970 0.0510 6.6270 0.9710 ;
      RECT 6.7490 0.0510 6.7790 0.9710 ;
      RECT 6.9010 0.0510 6.9310 0.9710 ;
      RECT 7.0530 0.0510 7.0830 0.9710 ;
      RECT 7.2050 0.0510 7.2350 0.9710 ;
      RECT 7.5090 0.0510 7.5390 0.9710 ;
      RECT 7.3570 0.0510 7.3870 0.9710 ;
      RECT 4.7730 2.3730 4.8030 3.2930 ;
      RECT 4.6210 2.3730 4.6510 3.2930 ;
      RECT 4.4690 2.3730 4.4990 3.2930 ;
      RECT 4.9250 2.3730 4.9550 3.2930 ;
      RECT 5.0770 2.3730 5.1070 3.2930 ;
      RECT 5.2290 2.3730 5.2590 3.2930 ;
      RECT 2.3410 2.3730 2.3710 3.2930 ;
      RECT 2.4930 2.3730 2.5230 3.2930 ;
      RECT 2.6450 2.3730 2.6750 3.2930 ;
      RECT 2.7970 2.3730 2.8270 3.2930 ;
      RECT 3.1010 2.3730 3.1310 3.2930 ;
      RECT 5.9890 0.0510 6.0190 1.9790 ;
      RECT 6.1410 0.0510 6.1710 1.9790 ;
      RECT 5.8370 0.0510 5.8670 1.9790 ;
      RECT 6.2930 0.0510 6.3230 1.9790 ;
      RECT 5.6850 0.0510 5.7150 0.9710 ;
      RECT 6.4450 0.0510 6.4750 0.9710 ;
      RECT 5.3810 1.3510 5.4110 2.1670 ;
      RECT 5.6850 1.3510 5.7150 1.9790 ;
      RECT 5.5330 1.3510 5.5630 1.9790 ;
      RECT 6.4450 1.3510 6.4750 1.9790 ;
      RECT 6.5970 1.3510 6.6270 1.9790 ;
      RECT 6.9010 1.3510 6.9310 1.8920 ;
      RECT 4.6210 0.0510 4.6510 1.9790 ;
      RECT 4.4690 0.0510 4.4990 1.9790 ;
      RECT 4.7730 0.0510 4.8030 1.9790 ;
      RECT 4.3170 0.0510 4.3470 1.9790 ;
      RECT 4.9250 0.0510 4.9550 0.9710 ;
      RECT 4.1650 0.0510 4.1950 0.9710 ;
      RECT 5.2290 1.3510 5.2590 2.1670 ;
      RECT 3.8610 1.3510 3.8910 2.1670 ;
      RECT 4.9250 1.3510 4.9550 1.9790 ;
      RECT 5.0770 1.3510 5.1070 1.9790 ;
      RECT 4.1650 1.3510 4.1950 1.9790 ;
      RECT 4.0130 1.3510 4.0430 1.9790 ;
      RECT 2.9490 0.0510 2.9790 1.9790 ;
      RECT 3.1010 0.0510 3.1310 1.9790 ;
      RECT 2.7970 0.0510 2.8270 1.9790 ;
      RECT 3.2530 0.0510 3.2830 1.9790 ;
    LAYER NWELL ;
      RECT -0.1150 2.3510 7.7150 3.4450 ;
      RECT 0.2310 1.8970 7.3680 2.3510 ;
      RECT 0.2310 1.0520 0.5940 1.8970 ;
      RECT 6.9650 1.0520 7.3680 1.8970 ;
      RECT 0.2310 0.9930 7.3680 1.0520 ;
      RECT -0.1150 -0.1010 7.7150 0.9930 ;
    LAYER M1 ;
      RECT 5.2000 1.9390 6.8400 1.9890 ;
      RECT 6.8150 1.7520 6.8650 1.9900 ;
      RECT 2.2550 1.7520 2.3050 1.9640 ;
      RECT 0.7600 1.9390 2.4000 1.9890 ;
      RECT 2.1600 1.9390 3.8000 1.9890 ;
      RECT 3.7750 1.7520 3.8250 1.9890 ;
      RECT 3.8000 1.9390 5.4400 1.9890 ;
      RECT 5.2950 1.7520 5.3450 1.9640 ;
      RECT 0.6690 1.9390 0.7840 1.9890 ;
      RECT 0.7350 1.7520 0.7850 1.9640 ;
      RECT 0.6690 2.2640 0.7850 2.3140 ;
      RECT 0.7350 2.2640 0.7850 3.2300 ;
      RECT 0.6690 1.9890 0.7190 2.2640 ;
  END
END FOOT2X16_LVT

MACRO FOOT2X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.128 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VSSG
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.7500 1.1750 0.9940 1.2570 ;
        RECT 0.8860 1.2570 0.9360 1.5330 ;
        RECT 0.8710 1.5330 1.5610 1.5890 ;
    END
  END VSSG

  PIN VSS
    DIRECTION OUTPUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.1280 1.7020 ;
        RECT 1.0390 1.7020 1.0890 1.8320 ;
    END
  END VSS

  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8060 2.0730 0.9820 2.1830 ;
    END
    ANTENNAGATEAREA 0.0366 ;
  END SLEEP

  PIN SLEEPOUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3130 1.1610 1.4230 1.2710 ;
        RECT 1.3430 1.2710 1.3930 1.4830 ;
        RECT 1.3430 0.1820 1.3930 1.1610 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END SLEEPOUT

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.1280 0.0300 ;
        RECT 1.4950 0.0300 1.5450 0.9290 ;
        RECT 1.1910 0.0300 1.2410 0.9290 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 2.1280 3.3740 ;
        RECT 0.8870 2.4400 0.9370 3.3140 ;
    END
  END VDD
  OBS
    LAYER NWELL ;
      RECT -0.1150 2.3510 2.2430 3.4450 ;
      RECT 0.2310 1.8970 1.8970 2.3510 ;
      RECT 0.2310 1.0520 0.6540 1.8970 ;
      RECT 1.6260 1.0520 1.8970 1.8970 ;
      RECT 0.2310 0.9930 1.8970 1.0520 ;
      RECT -0.1150 -0.1010 2.2430 0.9930 ;
    LAYER M1 ;
      RECT 0.7600 1.9390 1.4850 1.9890 ;
      RECT 0.6690 1.9390 0.7840 1.9890 ;
      RECT 0.7350 1.7570 0.7850 1.9710 ;
      RECT 0.6690 2.2640 0.7850 2.3140 ;
      RECT 0.7350 2.2640 0.7850 3.2300 ;
      RECT 0.6690 1.9890 0.7190 2.2640 ;
    LAYER PO ;
      RECT 0.5170 2.3730 0.5470 3.2930 ;
      RECT 0.3650 2.3730 0.3950 3.2930 ;
      RECT 0.2130 2.3730 0.2430 3.2930 ;
      RECT 0.0610 2.3730 0.0910 3.2930 ;
      RECT 0.5170 1.3510 0.5470 1.8920 ;
      RECT 0.3650 1.3510 0.3950 1.8920 ;
      RECT 0.2130 1.3510 0.2430 1.8920 ;
      RECT 0.0610 1.3510 0.0910 1.8920 ;
      RECT 0.9730 0.0510 1.0030 0.9710 ;
      RECT 0.8210 0.0510 0.8510 0.9710 ;
      RECT 0.3650 0.0510 0.3950 0.9710 ;
      RECT 0.2130 0.0510 0.2430 0.9710 ;
      RECT 0.0610 0.0510 0.0910 0.9710 ;
      RECT 0.6690 0.0510 0.6990 0.9710 ;
      RECT 0.5170 0.0510 0.5470 0.9710 ;
      RECT 2.0370 1.3510 2.0670 1.8920 ;
      RECT 1.7330 0.0510 1.7630 0.9710 ;
      RECT 1.5810 0.0510 1.6110 0.9710 ;
      RECT 2.0370 0.0510 2.0670 0.9710 ;
      RECT 1.8850 0.0510 1.9150 0.9710 ;
      RECT 1.8850 1.3510 1.9150 1.8920 ;
      RECT 1.7330 1.3510 1.7630 1.8920 ;
      RECT 2.0370 2.3730 2.0670 3.2930 ;
      RECT 1.8850 2.3730 1.9150 3.2930 ;
      RECT 1.7330 2.3730 1.7630 3.2930 ;
      RECT 1.5810 2.3730 1.6110 3.2930 ;
      RECT 1.4290 2.3730 1.4590 3.2930 ;
      RECT 1.1250 2.3730 1.1550 3.2930 ;
      RECT 1.2770 2.3730 1.3070 3.2930 ;
      RECT 0.9730 2.3730 1.0030 3.2930 ;
      RECT 1.4290 0.0510 1.4590 1.9790 ;
      RECT 1.1250 0.0510 1.1550 0.9710 ;
      RECT 0.6690 2.3730 0.6990 3.2930 ;
      RECT 1.2770 0.0510 1.3070 1.9790 ;
      RECT 0.6690 1.3510 0.6990 1.8920 ;
      RECT 0.8210 1.3510 0.8510 3.2930 ;
      RECT 1.1250 1.3510 1.1550 1.9790 ;
      RECT 0.9730 1.3510 1.0030 1.9790 ;
      RECT 1.5810 1.3510 1.6110 1.9630 ;
  END
END FOOT2X2_LVT

MACRO FOOT2X32_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 13.68 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VSSG
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.7500 1.1750 0.9940 1.2570 ;
        RECT 0.8860 1.2570 0.9360 1.5350 ;
        RECT 0.8710 1.5350 12.8090 1.5910 ;
    END
  END VSSG

  PIN VSS
    DIRECTION OUTPUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 13.6800 1.7020 ;
        RECT 4.9910 1.7020 5.0410 1.8320 ;
        RECT 4.0790 1.7020 4.1290 1.8320 ;
        RECT 2.5590 1.7020 2.6090 1.8320 ;
        RECT 3.4710 1.7020 3.5210 1.8320 ;
        RECT 1.9510 1.7020 2.0010 1.8320 ;
        RECT 1.0390 1.7020 1.0890 1.8320 ;
        RECT 8.0310 1.7020 8.0810 1.8320 ;
        RECT 7.1190 1.7020 7.1690 1.8320 ;
        RECT 8.6390 1.7020 8.6890 1.8320 ;
        RECT 9.5510 1.7020 9.6010 1.8320 ;
        RECT 11.0710 1.7020 11.1210 1.8320 ;
        RECT 10.1590 1.7020 10.2090 1.8320 ;
        RECT 11.6790 1.7020 11.7290 1.8320 ;
        RECT 12.5910 1.7020 12.6410 1.8320 ;
        RECT 5.5990 1.7020 5.6490 1.8320 ;
        RECT 6.5110 1.7020 6.5610 1.8320 ;
    END
  END VSS

  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8000 2.1560 0.9670 2.1830 ;
        RECT 0.8000 2.1060 12.9180 2.1560 ;
        RECT 0.8000 2.0730 0.9670 2.1060 ;
    END
    ANTENNAGATEAREA 0.2256 ;
  END SLEEP

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 13.6800 0.0300 ;
        RECT 2.7110 0.0300 2.7610 0.9240 ;
        RECT 3.0150 0.0300 3.0650 0.9240 ;
        RECT 3.3190 0.0300 3.3690 0.9240 ;
        RECT 1.7990 0.0300 1.8490 0.9240 ;
        RECT 1.4950 0.0300 1.5450 0.9240 ;
        RECT 1.1910 0.0300 1.2410 0.9240 ;
        RECT 10.9190 0.0300 10.9690 0.9240 ;
        RECT 10.6150 0.0300 10.6650 0.9240 ;
        RECT 11.8310 0.0300 11.8810 0.9240 ;
        RECT 12.1350 0.0300 12.1850 0.9240 ;
        RECT 12.4390 0.0300 12.4890 0.9240 ;
        RECT 7.8790 0.0300 7.9290 0.9240 ;
        RECT 7.5750 0.0300 7.6250 0.9240 ;
        RECT 7.2710 0.0300 7.3210 0.9240 ;
        RECT 8.7910 0.0300 8.8410 0.9240 ;
        RECT 9.0950 0.0300 9.1450 0.9240 ;
        RECT 9.3990 0.0300 9.4490 0.9240 ;
        RECT 10.3110 0.0300 10.3610 0.9240 ;
        RECT 5.7510 0.0300 5.8010 0.9240 ;
        RECT 6.0550 0.0300 6.1050 0.9240 ;
        RECT 6.3590 0.0300 6.4090 0.9240 ;
        RECT 4.8390 0.0300 4.8890 0.9240 ;
        RECT 4.5350 0.0300 4.5850 0.9240 ;
        RECT 4.2310 0.0300 4.2810 0.9240 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 13.6800 3.3740 ;
        RECT 0.8870 2.4890 0.9370 3.3140 ;
    END
  END VDD

  PIN SLEEPOUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 12.2870 1.2710 12.3370 1.4840 ;
        RECT 11.9830 1.2000 12.0330 1.4840 ;
        RECT 10.4630 1.2000 10.5130 1.4840 ;
        RECT 10.7670 1.2000 10.8170 1.4840 ;
        RECT 9.2470 1.2000 9.2970 1.4840 ;
        RECT 8.9430 1.2000 8.9930 1.4840 ;
        RECT 7.4230 1.2000 7.4730 1.4840 ;
        RECT 7.7270 1.2000 7.7770 1.4840 ;
        RECT 12.2570 1.2000 12.3670 1.2710 ;
        RECT 6.2070 1.2000 6.2570 1.4840 ;
        RECT 5.9030 1.2000 5.9530 1.4840 ;
        RECT 4.6870 1.2000 4.7370 1.4840 ;
        RECT 3.1670 1.2000 3.2170 1.4840 ;
        RECT 4.3830 1.2000 4.4330 1.4840 ;
        RECT 1.6470 1.2000 1.6970 1.4840 ;
        RECT 2.8630 1.2000 2.9130 1.4840 ;
        RECT 1.3430 1.2000 1.3930 1.4840 ;
        RECT 1.3430 1.1610 12.3670 1.2000 ;
        RECT 1.3430 1.1500 12.3370 1.1610 ;
        RECT 12.2870 0.1980 12.3370 1.1500 ;
        RECT 11.9830 0.1980 12.0330 1.1500 ;
        RECT 10.4630 0.1980 10.5130 1.1500 ;
        RECT 10.7670 0.1980 10.8170 1.1500 ;
        RECT 9.2470 0.1980 9.2970 1.1500 ;
        RECT 8.9430 0.1980 8.9930 1.1500 ;
        RECT 7.4230 0.1980 7.4730 1.1500 ;
        RECT 7.7270 0.1980 7.7770 1.1500 ;
        RECT 6.2070 0.1980 6.2570 1.1500 ;
        RECT 5.9030 0.1980 5.9530 1.1500 ;
        RECT 4.6870 0.1980 4.7370 1.1500 ;
        RECT 3.1670 0.1980 3.2170 1.1500 ;
        RECT 4.3830 0.1980 4.4330 1.1500 ;
        RECT 1.6470 0.1980 1.6970 1.1500 ;
        RECT 2.8630 0.1980 2.9130 1.1500 ;
        RECT 1.3430 0.1980 1.3930 1.1500 ;
    END
    ANTENNADIFFAREA 2.3808 ;
  END SLEEPOUT
  OBS
    LAYER PO ;
      RECT 13.4370 2.3730 13.4670 3.2930 ;
      RECT 13.5890 2.3730 13.6190 3.2930 ;
      RECT 13.2850 2.3730 13.3150 3.2930 ;
      RECT 12.8290 2.3730 12.8590 3.2930 ;
      RECT 12.9810 2.3730 13.0110 3.2930 ;
      RECT 12.6770 2.3730 12.7070 3.2930 ;
      RECT 13.5890 1.3510 13.6190 1.8920 ;
      RECT 13.4370 1.3510 13.4670 1.8920 ;
      RECT 13.2850 1.3510 13.3150 1.8920 ;
      RECT 13.1330 1.3510 13.1630 1.8920 ;
      RECT 5.8370 0.0510 5.8670 1.9790 ;
      RECT 6.2930 0.0510 6.3230 1.9790 ;
      RECT 5.6850 0.0510 5.7150 0.9710 ;
      RECT 6.4450 0.0510 6.4750 0.9710 ;
      RECT 5.6850 1.3510 5.7150 1.9790 ;
      RECT 6.4450 1.3510 6.4750 1.9790 ;
      RECT 6.5970 1.3510 6.6270 1.9790 ;
      RECT 6.5970 0.0510 6.6270 0.9710 ;
      RECT 6.4450 2.3730 6.4750 3.2930 ;
      RECT 6.5970 2.3730 6.6270 3.2930 ;
      RECT 5.6850 2.3730 5.7150 3.2930 ;
      RECT 5.8370 2.3730 5.8670 3.2930 ;
      RECT 6.1410 2.3730 6.1710 3.2930 ;
      RECT 6.2930 2.3730 6.3230 3.2930 ;
      RECT 5.9890 2.3730 6.0190 3.2930 ;
      RECT 6.9010 2.3730 6.9310 3.2930 ;
      RECT 7.6610 0.0510 7.6910 1.9790 ;
      RECT 7.5090 0.0510 7.5390 1.9790 ;
      RECT 7.3570 0.0510 7.3870 1.9790 ;
      RECT 7.2050 0.0510 7.2350 0.9710 ;
      RECT 6.9010 1.3510 6.9310 2.1670 ;
      RECT 7.2050 1.3510 7.2350 1.9790 ;
      RECT 7.0530 1.3510 7.0830 1.9790 ;
      RECT 6.7490 1.3510 6.7790 2.1670 ;
      RECT 7.0530 0.0510 7.0830 0.9710 ;
      RECT 6.9010 0.0510 6.9310 0.9710 ;
      RECT 6.7490 0.0510 6.7790 0.9710 ;
      RECT 7.6610 2.3730 7.6910 3.2930 ;
      RECT 7.0530 2.3730 7.0830 3.2930 ;
      RECT 7.3570 2.3730 7.3870 3.2930 ;
      RECT 7.5090 2.3730 7.5390 3.2930 ;
      RECT 7.2050 2.3730 7.2350 3.2930 ;
      RECT 6.7490 2.3730 6.7790 3.2930 ;
      RECT 8.5730 1.3510 8.6030 1.9790 ;
      RECT 7.8130 0.0510 7.8430 1.9790 ;
      RECT 7.9650 0.0510 7.9950 0.9710 ;
      RECT 8.2690 1.3510 8.2990 2.1670 ;
      RECT 7.9650 1.3510 7.9950 1.9790 ;
      RECT 8.1170 1.3510 8.1470 1.9790 ;
      RECT 8.4210 0.0510 8.4510 0.9710 ;
      RECT 8.2690 0.0510 8.2990 0.9710 ;
      RECT 8.5730 0.0510 8.6030 0.9710 ;
      RECT 8.1170 0.0510 8.1470 0.9710 ;
      RECT 8.4210 1.3510 8.4510 2.1670 ;
      RECT 8.1170 2.3730 8.1470 3.2930 ;
      RECT 7.9650 2.3730 7.9950 3.2930 ;
      RECT 8.4210 2.3730 8.4510 3.2930 ;
      RECT 8.5730 2.3730 8.6030 3.2930 ;
      RECT 8.2690 2.3730 8.2990 3.2930 ;
      RECT 7.8130 2.3730 7.8430 3.2930 ;
      RECT 8.7250 1.3510 8.7550 1.9790 ;
      RECT 9.4850 1.3510 9.5150 1.9790 ;
      RECT 9.6370 1.3510 9.6670 1.9790 ;
      RECT 9.0290 0.0510 9.0590 1.9790 ;
      RECT 9.1810 0.0510 9.2110 1.9790 ;
      RECT 9.6370 0.0510 9.6670 0.9710 ;
      RECT 8.8770 0.0510 8.9070 1.9790 ;
      RECT 9.3330 0.0510 9.3630 1.9790 ;
      RECT 8.7250 0.0510 8.7550 0.9710 ;
      RECT 9.4850 0.0510 9.5150 0.9710 ;
      RECT 8.7250 2.3730 8.7550 3.2930 ;
      RECT 9.0290 2.3730 9.0590 3.2930 ;
      RECT 9.3330 2.3730 9.3630 3.2930 ;
      RECT 9.1810 2.3730 9.2110 3.2930 ;
      RECT 9.6370 2.3730 9.6670 3.2930 ;
      RECT 9.4850 2.3730 9.5150 3.2930 ;
      RECT 8.8770 2.3730 8.9070 3.2930 ;
      RECT 9.7890 0.0510 9.8190 0.9710 ;
      RECT 9.9410 0.0510 9.9710 0.9710 ;
      RECT 10.0930 0.0510 10.1230 0.9710 ;
      RECT 10.5490 0.0510 10.5790 1.9790 ;
      RECT 10.3970 0.0510 10.4270 1.9790 ;
      RECT 10.2450 0.0510 10.2750 0.9710 ;
      RECT 10.2450 1.3510 10.2750 1.9790 ;
      RECT 10.0930 1.3510 10.1230 1.9790 ;
      RECT 9.7890 1.3510 9.8190 2.1670 ;
      RECT 9.9410 1.3510 9.9710 2.1670 ;
      RECT 9.7890 2.3730 9.8190 3.2930 ;
      RECT 9.9410 2.3730 9.9710 3.2930 ;
      RECT 10.0930 2.3730 10.1230 3.2930 ;
      RECT 10.3970 2.3730 10.4270 3.2930 ;
      RECT 10.5490 2.3730 10.5790 3.2930 ;
      RECT 10.2450 2.3730 10.2750 3.2930 ;
      RECT 11.1570 0.0510 11.1870 0.9710 ;
      RECT 11.6130 0.0510 11.6430 0.9710 ;
      RECT 11.3090 0.0510 11.3390 0.9710 ;
      RECT 11.4610 0.0510 11.4910 0.9710 ;
      RECT 11.6130 1.3510 11.6430 1.9790 ;
      RECT 10.7010 0.0510 10.7310 1.9790 ;
      RECT 10.8530 0.0510 10.8830 1.9790 ;
      RECT 11.0050 0.0510 11.0350 0.9710 ;
      RECT 11.3090 1.3510 11.3390 2.1670 ;
      RECT 11.4610 1.3510 11.4910 2.1670 ;
      RECT 11.0050 1.3510 11.0350 1.9790 ;
      RECT 11.1570 1.3510 11.1870 1.9790 ;
      RECT 10.7010 2.3730 10.7310 3.2930 ;
      RECT 11.0050 2.3730 11.0350 3.2930 ;
      RECT 11.1570 2.3730 11.1870 3.2930 ;
      RECT 10.8530 2.3730 10.8830 3.2930 ;
      RECT 11.4610 2.3730 11.4910 3.2930 ;
      RECT 11.6130 2.3730 11.6430 3.2930 ;
      RECT 11.3090 2.3730 11.3390 3.2930 ;
      RECT 12.0690 0.0510 12.0990 1.9790 ;
      RECT 12.2210 0.0510 12.2510 1.9790 ;
      RECT 11.9170 0.0510 11.9470 1.9790 ;
      RECT 12.3730 0.0510 12.4030 1.9790 ;
      RECT 11.7650 0.0510 11.7950 0.9710 ;
      RECT 12.5250 0.0510 12.5550 0.9710 ;
      RECT 11.7650 1.3510 11.7950 1.9790 ;
      RECT 12.5250 1.3510 12.5550 1.9790 ;
      RECT 11.7650 2.3730 11.7950 3.2930 ;
      RECT 12.0690 2.3730 12.0990 3.2930 ;
      RECT 12.3730 2.3730 12.4030 3.2930 ;
      RECT 12.2210 2.3730 12.2510 3.2930 ;
      RECT 11.9170 2.3730 11.9470 3.2930 ;
      RECT 12.5250 2.3730 12.5550 3.2930 ;
      RECT 12.8290 1.3510 12.8590 2.1670 ;
      RECT 12.8290 0.0510 12.8590 0.9710 ;
      RECT 12.6770 0.0510 12.7070 0.9710 ;
      RECT 13.5890 0.0510 13.6190 0.9710 ;
      RECT 13.4370 0.0510 13.4670 0.9710 ;
      RECT 13.2850 0.0510 13.3150 0.9710 ;
      RECT 13.1330 0.0510 13.1630 0.9710 ;
      RECT 12.9810 0.0510 13.0110 0.9710 ;
      RECT 12.6770 1.3510 12.7070 1.9790 ;
      RECT 12.9810 1.3510 13.0110 1.8920 ;
      RECT 13.1330 2.3730 13.1630 3.2930 ;
      RECT 0.6690 2.3730 0.6990 3.2930 ;
      RECT 0.6690 1.3510 0.6990 1.8920 ;
      RECT 0.5170 1.3510 0.5470 1.8920 ;
      RECT 0.3650 1.3510 0.3950 1.8920 ;
      RECT 0.2130 1.3510 0.2430 1.8920 ;
      RECT 0.0610 1.3510 0.0910 1.8920 ;
      RECT 0.5170 0.0510 0.5470 0.9710 ;
      RECT 0.2130 0.0510 0.2430 0.9710 ;
      RECT 0.3650 0.0510 0.3950 0.9710 ;
      RECT 0.0610 0.0510 0.0910 0.9710 ;
      RECT 0.6690 0.0510 0.6990 0.9710 ;
      RECT 0.0610 2.3730 0.0910 3.2930 ;
      RECT 0.3650 2.3730 0.3950 3.2930 ;
      RECT 0.5170 2.3730 0.5470 3.2930 ;
      RECT 0.2130 2.3730 0.2430 3.2930 ;
      RECT 1.5810 0.0510 1.6110 1.9790 ;
      RECT 0.9730 2.3730 1.0030 3.2930 ;
      RECT 1.4290 0.0510 1.4590 1.9790 ;
      RECT 1.1250 0.0510 1.1550 0.9710 ;
      RECT 1.2770 0.0510 1.3070 1.9790 ;
      RECT 0.8210 1.3510 0.8510 3.2930 ;
      RECT 1.1250 1.3510 1.1550 1.9790 ;
      RECT 0.9730 1.3510 1.0030 1.9790 ;
      RECT 1.5810 2.3730 1.6110 3.2930 ;
      RECT 1.2770 2.3730 1.3070 3.2930 ;
      RECT 1.4290 2.3730 1.4590 3.2930 ;
      RECT 1.1250 2.3730 1.1550 3.2930 ;
      RECT 0.9730 0.0510 1.0030 0.9710 ;
      RECT 0.8210 0.0510 0.8510 0.9710 ;
      RECT 2.0370 1.3510 2.0670 1.9790 ;
      RECT 2.1890 1.3510 2.2190 2.1670 ;
      RECT 2.6450 0.0510 2.6750 0.9710 ;
      RECT 2.3410 1.3510 2.3710 2.1670 ;
      RECT 2.6450 1.3510 2.6750 1.9790 ;
      RECT 2.4930 1.3510 2.5230 1.9790 ;
      RECT 2.1890 0.0510 2.2190 0.9710 ;
      RECT 2.4930 0.0510 2.5230 0.9710 ;
      RECT 1.8850 2.3730 1.9150 3.2930 ;
      RECT 2.0370 2.3730 2.0670 3.2930 ;
      RECT 1.7330 2.3730 1.7630 3.2930 ;
      RECT 2.0370 0.0510 2.0670 0.9710 ;
      RECT 2.3410 0.0510 2.3710 0.9710 ;
      RECT 2.1890 2.3730 2.2190 3.2930 ;
      RECT 2.4930 2.3730 2.5230 3.2930 ;
      RECT 2.6450 2.3730 2.6750 3.2930 ;
      RECT 2.3410 2.3730 2.3710 3.2930 ;
      RECT 1.7330 0.0510 1.7630 1.9790 ;
      RECT 1.8850 0.0510 1.9150 0.9710 ;
      RECT 1.8850 1.3510 1.9150 1.9790 ;
      RECT 2.9490 0.0510 2.9790 1.9790 ;
      RECT 3.1010 0.0510 3.1310 1.9790 ;
      RECT 2.7970 0.0510 2.8270 1.9790 ;
      RECT 3.2530 0.0510 3.2830 1.9790 ;
      RECT 3.4050 0.0510 3.4350 0.9710 ;
      RECT 3.4050 1.3510 3.4350 1.9790 ;
      RECT 3.5570 1.3510 3.5870 1.9790 ;
      RECT 3.5570 0.0510 3.5870 0.9710 ;
      RECT 3.5570 2.3730 3.5870 3.2930 ;
      RECT 3.4050 2.3730 3.4350 3.2930 ;
      RECT 3.2530 2.3730 3.2830 3.2930 ;
      RECT 2.7970 2.3730 2.8270 3.2930 ;
      RECT 3.1010 2.3730 3.1310 3.2930 ;
      RECT 2.9490 2.3730 2.9790 3.2930 ;
      RECT 3.7090 1.3510 3.7390 2.1670 ;
      RECT 4.6210 0.0510 4.6510 1.9790 ;
      RECT 4.4690 0.0510 4.4990 1.9790 ;
      RECT 4.3170 0.0510 4.3470 1.9790 ;
      RECT 4.1650 0.0510 4.1950 0.9710 ;
      RECT 3.8610 1.3510 3.8910 2.1670 ;
      RECT 4.1650 1.3510 4.1950 1.9790 ;
      RECT 4.0130 1.3510 4.0430 1.9790 ;
      RECT 3.7090 0.0510 3.7390 0.9710 ;
      RECT 3.8610 0.0510 3.8910 0.9710 ;
      RECT 4.0130 0.0510 4.0430 0.9710 ;
      RECT 4.6210 2.3730 4.6510 3.2930 ;
      RECT 3.8610 2.3730 3.8910 3.2930 ;
      RECT 3.7090 2.3730 3.7390 3.2930 ;
      RECT 4.1650 2.3730 4.1950 3.2930 ;
      RECT 4.4690 2.3730 4.4990 3.2930 ;
      RECT 4.3170 2.3730 4.3470 3.2930 ;
      RECT 4.0130 2.3730 4.0430 3.2930 ;
      RECT 5.3810 1.3510 5.4110 2.1670 ;
      RECT 5.5330 1.3510 5.5630 1.9790 ;
      RECT 4.7730 0.0510 4.8030 1.9790 ;
      RECT 4.9250 0.0510 4.9550 0.9710 ;
      RECT 5.2290 1.3510 5.2590 2.1670 ;
      RECT 4.9250 1.3510 4.9550 1.9790 ;
      RECT 5.0770 1.3510 5.1070 1.9790 ;
      RECT 5.5330 0.0510 5.5630 0.9710 ;
      RECT 5.2290 0.0510 5.2590 0.9710 ;
      RECT 5.3810 0.0510 5.4110 0.9710 ;
      RECT 5.0770 0.0510 5.1070 0.9710 ;
      RECT 4.7730 2.3730 4.8030 3.2930 ;
      RECT 5.0770 2.3730 5.1070 3.2930 ;
      RECT 4.9250 2.3730 4.9550 3.2930 ;
      RECT 5.3810 2.3730 5.4110 3.2930 ;
      RECT 5.5330 2.3730 5.5630 3.2930 ;
      RECT 5.2290 2.3730 5.2590 3.2930 ;
      RECT 5.9890 0.0510 6.0190 1.9790 ;
      RECT 6.1410 0.0510 6.1710 1.9790 ;
    LAYER NWELL ;
      RECT -0.0700 2.3510 13.7500 3.4450 ;
      RECT 0.2920 1.8970 13.4660 2.3510 ;
      RECT 0.2920 1.0520 0.6540 1.8970 ;
      RECT 13.0650 1.0520 13.4660 1.8970 ;
      RECT 0.2920 0.9930 13.4660 1.0520 ;
      RECT -0.0700 -0.1010 13.7500 0.9930 ;
    LAYER M1 ;
      RECT 11.2800 1.9390 12.9200 1.9890 ;
      RECT 12.8950 1.7520 12.9450 1.9910 ;
      RECT 2.2550 1.7520 2.3050 1.9640 ;
      RECT 0.7600 1.9390 2.4000 1.9890 ;
      RECT 2.1600 1.9390 3.8000 1.9890 ;
      RECT 3.7750 1.7520 3.8250 1.9890 ;
      RECT 3.8000 1.9390 5.4400 1.9890 ;
      RECT 5.2950 1.7520 5.3450 1.9640 ;
      RECT 5.2000 1.9390 6.8400 1.9890 ;
      RECT 6.8150 1.7520 6.8650 1.9900 ;
      RECT 6.8400 1.9390 8.4800 1.9890 ;
      RECT 8.3350 1.7520 8.3850 1.9640 ;
      RECT 8.2400 1.9390 9.8800 1.9890 ;
      RECT 9.8550 1.7520 9.9050 1.9890 ;
      RECT 9.8800 1.9390 11.5200 1.9890 ;
      RECT 11.3750 1.7520 11.4250 1.9640 ;
      RECT 0.6690 1.9390 0.7840 1.9890 ;
      RECT 0.7350 1.7520 0.7850 1.9640 ;
      RECT 0.6690 2.2640 0.7850 2.3140 ;
      RECT 0.7350 2.2640 0.7850 3.2150 ;
      RECT 0.6690 1.9890 0.7190 2.2640 ;
  END
END FOOT2X32_LVT

MACRO FOOT2X4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.192 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SLEEPOUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6470 1.2710 1.6970 1.4830 ;
        RECT 1.6170 1.2000 1.7270 1.2710 ;
        RECT 1.3430 1.1610 1.7270 1.2000 ;
        RECT 1.3430 1.1500 1.6970 1.1610 ;
        RECT 1.3430 1.2000 1.3930 1.4830 ;
        RECT 1.3430 0.1980 1.3930 1.1500 ;
        RECT 1.6470 0.1980 1.6970 1.1500 ;
    END
    ANTENNADIFFAREA 0.2976 ;
  END SLEEPOUT

  PIN VSSG
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.6910 1.1750 0.9360 1.2570 ;
        RECT 0.8860 1.2570 0.9360 1.5330 ;
        RECT 0.8710 1.5330 2.1880 1.5890 ;
    END
  END VSSG

  PIN VSS
    DIRECTION OUTPUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.1920 1.7020 ;
        RECT 1.9510 1.7020 2.0010 1.8320 ;
        RECT 1.0390 1.7020 1.0890 1.8320 ;
    END
  END VSS

  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7990 2.0730 0.9770 2.1060 ;
        RECT 0.7990 2.1060 2.2450 2.1560 ;
        RECT 0.7990 2.1560 0.9770 2.1830 ;
    END
    ANTENNAGATEAREA 0.0492 ;
  END SLEEP

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.1920 0.0300 ;
        RECT 1.7990 0.0300 1.8490 0.9240 ;
        RECT 1.4950 0.0300 1.5450 0.9240 ;
        RECT 1.1910 0.0300 1.2410 0.9240 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 3.1920 3.3740 ;
        RECT 0.8870 2.4880 0.9370 3.3140 ;
    END
  END VDD
  OBS
    LAYER NWELL ;
      RECT -0.1150 2.3510 3.3070 3.4450 ;
      RECT 0.2310 1.8970 2.9610 2.3510 ;
      RECT 0.2310 1.0520 0.5940 1.8970 ;
      RECT 2.5640 1.0520 2.9610 1.8970 ;
      RECT 0.2310 0.9930 2.9610 1.0520 ;
      RECT -0.1150 -0.1010 3.3070 0.9930 ;
    LAYER M1 ;
      RECT 2.2550 1.7520 2.3050 1.9640 ;
      RECT 0.7600 1.9390 2.4000 1.9890 ;
      RECT 0.6690 1.9390 0.7840 1.9890 ;
      RECT 0.7350 1.7540 0.7850 1.9640 ;
      RECT 0.6690 2.2640 0.7850 2.3140 ;
      RECT 0.7350 2.2640 0.7850 3.2140 ;
      RECT 0.6690 1.9890 0.7190 2.2640 ;
    LAYER PO ;
      RECT 2.9490 0.0510 2.9790 0.9710 ;
      RECT 2.7970 0.0510 2.8270 0.9710 ;
      RECT 2.6450 0.0510 2.6750 0.9710 ;
      RECT 2.3410 0.0510 2.3710 0.9710 ;
      RECT 2.7970 2.3730 2.8270 3.2930 ;
      RECT 0.9730 2.3730 1.0030 3.2930 ;
      RECT 1.4290 0.0510 1.4590 1.9790 ;
      RECT 1.1250 0.0510 1.1550 0.9710 ;
      RECT 0.6690 2.3730 0.6990 3.2930 ;
      RECT 1.2770 0.0510 1.3070 1.9790 ;
      RECT 0.6690 1.3510 0.6990 2.1670 ;
      RECT 2.1890 0.0510 2.2190 0.9710 ;
      RECT 0.8210 1.3510 0.8510 3.2930 ;
      RECT 1.1250 1.3510 1.1550 1.9790 ;
      RECT 0.9730 1.3510 1.0030 1.9790 ;
      RECT 2.0370 0.0510 2.0670 0.9710 ;
      RECT 0.0610 1.3510 0.0910 2.1670 ;
      RECT 0.5170 1.3510 0.5470 2.1670 ;
      RECT 0.3650 1.3510 0.3950 2.1670 ;
      RECT 0.2130 1.3510 0.2430 2.1670 ;
      RECT 1.8850 2.3730 1.9150 3.2930 ;
      RECT 2.1890 2.3730 2.2190 3.2930 ;
      RECT 2.3410 2.3730 2.3710 3.2930 ;
      RECT 2.0370 2.3730 2.0670 3.2930 ;
      RECT 1.1250 2.3730 1.1550 3.2930 ;
      RECT 1.4290 2.3730 1.4590 3.2930 ;
      RECT 2.9490 2.3730 2.9790 3.2930 ;
      RECT 1.5810 0.0510 1.6110 1.9790 ;
      RECT 1.7330 0.0510 1.7630 1.9790 ;
      RECT 0.2130 2.3730 0.2430 3.2930 ;
      RECT 1.8850 0.0510 1.9150 0.9710 ;
      RECT 1.8850 1.3510 1.9150 1.9790 ;
      RECT 2.0370 1.3510 2.0670 1.9790 ;
      RECT 2.4930 2.3730 2.5230 3.2930 ;
      RECT 2.6450 2.3730 2.6750 3.2930 ;
      RECT 0.5170 0.0510 0.5470 0.9710 ;
      RECT 0.0610 2.3730 0.0910 3.2930 ;
      RECT 1.7330 2.3730 1.7630 3.2930 ;
      RECT 0.3650 2.3730 0.3950 3.2930 ;
      RECT 1.5810 2.3730 1.6110 3.2930 ;
      RECT 1.2770 2.3730 1.3070 3.2930 ;
      RECT 3.1010 2.3730 3.1310 3.2930 ;
      RECT 0.5170 2.3730 0.5470 3.2930 ;
      RECT 2.3410 1.3510 2.3710 2.1670 ;
      RECT 0.9730 0.0510 1.0030 0.9710 ;
      RECT 0.8210 0.0510 0.8510 0.9710 ;
      RECT 0.6690 0.0510 0.6990 0.9710 ;
      RECT 2.1890 1.3510 2.2190 2.1670 ;
      RECT 0.3650 0.0510 0.3950 0.9710 ;
      RECT 0.2130 0.0510 0.2430 0.9710 ;
      RECT 0.0610 0.0510 0.0910 0.9710 ;
      RECT 3.1010 1.3510 3.1310 2.1670 ;
      RECT 2.9490 1.3510 2.9790 2.1670 ;
      RECT 2.7970 1.3510 2.8270 2.1670 ;
      RECT 2.6450 1.3510 2.6750 2.1670 ;
      RECT 2.4930 1.3510 2.5230 2.1670 ;
      RECT 2.4930 0.0510 2.5230 0.9710 ;
      RECT 3.1010 0.0510 3.1310 0.9710 ;
  END
END FOOT2X4_LVT

MACRO FOOT2X8_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.56 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SLEEPOUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.1370 1.2000 3.2470 1.2710 ;
        RECT 3.1670 1.2710 3.2170 1.4830 ;
        RECT 1.3430 1.1610 3.2470 1.2000 ;
        RECT 2.8630 1.2000 2.9130 1.4830 ;
        RECT 1.6470 1.2000 1.6970 1.4830 ;
        RECT 1.3430 1.2000 1.3930 1.4830 ;
        RECT 1.3430 1.1500 3.2170 1.1610 ;
        RECT 3.1670 0.1980 3.2170 1.1500 ;
        RECT 2.8630 0.1980 2.9130 1.1500 ;
        RECT 1.6470 0.1980 1.6970 1.1500 ;
        RECT 1.3430 0.1980 1.3930 1.1500 ;
    END
    ANTENNADIFFAREA 0.5952 ;
  END SLEEPOUT

  PIN VSSG
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.7500 1.1750 0.9940 1.2570 ;
        RECT 0.8860 1.2570 0.9360 1.5330 ;
        RECT 0.8710 1.5330 3.6890 1.5890 ;
    END
  END VSSG

  PIN VSS
    DIRECTION OUTPUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.5600 1.7020 ;
        RECT 2.5590 1.7020 2.6090 1.8320 ;
        RECT 3.4710 1.7020 3.5210 1.8320 ;
        RECT 1.9510 1.7020 2.0010 1.8320 ;
        RECT 1.0390 1.7020 1.0890 1.8320 ;
    END
  END VSS

  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8120 2.0710 0.9670 2.1060 ;
        RECT 0.8120 2.1060 3.7710 2.1560 ;
        RECT 0.8120 2.1560 0.9670 2.1810 ;
    END
    ANTENNAGATEAREA 0.0744 ;
  END SLEEP

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.5600 0.0300 ;
        RECT 2.7110 0.0300 2.7610 0.9240 ;
        RECT 3.0150 0.0300 3.0650 0.9240 ;
        RECT 3.3190 0.0300 3.3690 0.9240 ;
        RECT 1.7990 0.0300 1.8490 0.9240 ;
        RECT 1.4950 0.0300 1.5450 0.9240 ;
        RECT 1.1910 0.0300 1.2410 0.9240 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 4.5600 3.3740 ;
        RECT 0.8870 2.4880 0.9370 3.3140 ;
    END
  END VDD
  OBS
    LAYER NWELL ;
      RECT -0.1100 2.3510 4.6300 3.4450 ;
      RECT 0.2330 1.8970 4.3290 2.3510 ;
      RECT 0.2330 1.0520 0.6010 1.8970 ;
      RECT 3.9100 1.0520 4.3290 1.8970 ;
      RECT 0.2330 0.9930 4.3290 1.0520 ;
      RECT -0.0990 -0.1010 4.6300 0.9930 ;
    LAYER M1 ;
      RECT 2.1600 1.9390 3.8000 1.9890 ;
      RECT 3.7750 1.7520 3.8250 1.9890 ;
      RECT 2.2550 1.7520 2.3050 1.9640 ;
      RECT 0.7600 1.9390 2.4000 1.9890 ;
      RECT 0.6690 1.9390 0.7840 1.9890 ;
      RECT 0.7350 1.7520 0.7850 1.9640 ;
      RECT 0.6690 2.2640 0.7850 2.3140 ;
      RECT 0.7350 2.2640 0.7850 3.2140 ;
      RECT 0.6690 1.9890 0.7190 2.2640 ;
    LAYER PO ;
      RECT 3.1010 0.0510 3.1310 1.9790 ;
      RECT 2.7970 0.0510 2.8270 1.9790 ;
      RECT 3.2530 0.0510 3.2830 1.9790 ;
      RECT 2.6450 0.0510 2.6750 0.9710 ;
      RECT 3.4050 0.0510 3.4350 0.9710 ;
      RECT 2.3410 1.3510 2.3710 2.1670 ;
      RECT 2.6450 1.3510 2.6750 1.9790 ;
      RECT 2.4930 1.3510 2.5230 1.9790 ;
      RECT 3.4050 1.3510 3.4350 1.9790 ;
      RECT 3.5570 1.3510 3.5870 1.9790 ;
      RECT 2.9490 0.0510 2.9790 1.9790 ;
      RECT 3.8610 1.3510 3.8910 1.8920 ;
      RECT 1.5810 0.0510 1.6110 1.9790 ;
      RECT 1.7330 0.0510 1.7630 1.9790 ;
      RECT 1.8850 0.0510 1.9150 0.9710 ;
      RECT 1.8850 1.3510 1.9150 1.9790 ;
      RECT 2.0370 1.3510 2.0670 1.9790 ;
      RECT 3.7090 1.3510 3.7390 2.1670 ;
      RECT 2.1890 1.3510 2.2190 2.1670 ;
      RECT 0.9730 2.3730 1.0030 3.2930 ;
      RECT 1.4290 0.0510 1.4590 1.9790 ;
      RECT 1.1250 0.0510 1.1550 0.9710 ;
      RECT 0.6690 2.3730 0.6990 3.2930 ;
      RECT 1.2770 0.0510 1.3070 1.9790 ;
      RECT 0.6690 1.3510 0.6990 1.8920 ;
      RECT 0.8210 1.3510 0.8510 3.2930 ;
      RECT 1.1250 1.3510 1.1550 1.9790 ;
      RECT 0.9730 1.3510 1.0030 1.9790 ;
      RECT 3.8610 2.3730 3.8910 3.2930 ;
      RECT 3.7090 2.3730 3.7390 3.2930 ;
      RECT 2.7970 2.3730 2.8270 3.2930 ;
      RECT 2.9490 2.3730 2.9790 3.2930 ;
      RECT 3.1010 2.3730 3.1310 3.2930 ;
      RECT 3.2530 2.3730 3.2830 3.2930 ;
      RECT 3.4050 2.3730 3.4350 3.2930 ;
      RECT 3.5570 2.3730 3.5870 3.2930 ;
      RECT 1.8850 2.3730 1.9150 3.2930 ;
      RECT 2.0370 2.3730 2.0670 3.2930 ;
      RECT 2.1890 2.3730 2.2190 3.2930 ;
      RECT 2.3410 2.3730 2.3710 3.2930 ;
      RECT 2.4930 2.3730 2.5230 3.2930 ;
      RECT 2.6450 2.3730 2.6750 3.2930 ;
      RECT 1.7330 2.3730 1.7630 3.2930 ;
      RECT 1.5810 2.3730 1.6110 3.2930 ;
      RECT 1.4290 2.3730 1.4590 3.2930 ;
      RECT 1.2770 2.3730 1.3070 3.2930 ;
      RECT 1.1250 2.3730 1.1550 3.2930 ;
      RECT 3.8610 0.0510 3.8910 0.9710 ;
      RECT 3.7090 0.0510 3.7390 0.9710 ;
      RECT 3.5570 0.0510 3.5870 0.9710 ;
      RECT 2.4930 0.0510 2.5230 0.9710 ;
      RECT 2.3410 0.0510 2.3710 0.9710 ;
      RECT 2.1890 0.0510 2.2190 0.9710 ;
      RECT 2.0370 0.0510 2.0670 0.9710 ;
      RECT 0.6690 0.0510 0.6990 0.9710 ;
      RECT 0.8210 0.0510 0.8510 0.9710 ;
      RECT 0.9730 0.0510 1.0030 0.9710 ;
      RECT 4.0130 0.0610 4.0430 3.2810 ;
      RECT 4.1650 0.0610 4.1950 3.2810 ;
      RECT 4.3170 0.0610 4.3470 3.2810 ;
      RECT 4.4690 0.0610 4.4990 3.2810 ;
      RECT 0.0610 0.0610 0.0910 3.2810 ;
      RECT 0.2130 0.0610 0.2430 3.2810 ;
      RECT 0.3650 0.0610 0.3950 3.2810 ;
      RECT 0.5170 0.0610 0.5470 3.2810 ;
  END
END FOOT2X8_LVT

MACRO DFFNARX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.408 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.4080 0.0300 ;
        RECT 0.5860 0.0300 0.6360 0.1960 ;
        RECT 0.2790 0.0300 0.3290 0.4190 ;
        RECT 3.7750 0.0300 3.8250 0.2200 ;
        RECT 3.4710 0.0300 3.5210 0.3300 ;
        RECT 1.5410 0.0300 1.5910 0.2870 ;
        RECT 0.5860 0.1960 0.9370 0.2460 ;
        RECT 2.9990 0.3300 3.5370 0.3800 ;
        RECT 1.5410 0.2870 2.0010 0.3370 ;
        RECT 0.8870 0.2460 0.9370 0.4500 ;
        RECT 0.7350 0.2460 0.7850 0.4500 ;
        RECT 1.9510 0.3370 2.0010 0.4610 ;
        RECT 1.9510 0.2490 2.0010 0.2870 ;
        RECT 1.9510 0.1990 2.1760 0.2490 ;
    END
  END VSS

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0490 1.1610 4.1600 1.2210 ;
        RECT 3.9270 1.2210 4.1600 1.2710 ;
        RECT 4.1090 0.2040 4.1590 1.1610 ;
        RECT 3.9270 1.2710 3.9770 1.5460 ;
        RECT 3.9110 0.1540 4.1590 0.2040 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.4080 1.7020 ;
        RECT 0.2790 1.0330 0.3290 1.6420 ;
        RECT 3.7750 0.9470 3.8250 1.6420 ;
        RECT 2.1270 1.3280 2.1770 1.6420 ;
        RECT 3.5110 1.3580 3.5610 1.6420 ;
        RECT 0.4330 1.3640 0.4830 1.6420 ;
        RECT 1.9340 1.2780 2.1770 1.3280 ;
        RECT 2.8340 1.3080 3.5610 1.3580 ;
        RECT 0.4330 1.3440 0.9370 1.3640 ;
        RECT 0.4340 1.3140 0.9370 1.3440 ;
        RECT 0.7350 1.0980 0.7850 1.3140 ;
        RECT 0.8870 1.1110 0.9370 1.3140 ;
    END
  END VDD

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7230 0.0890 2.8530 0.1390 ;
        RECT 2.7710 0.1390 2.8530 0.1750 ;
        RECT 1.7230 0.1390 1.8790 0.2070 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.3590 0.6800 ;
        RECT 0.2490 0.6800 0.4210 0.7300 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.4240 0.7250 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8970 1.0090 4.0070 1.1190 ;
        RECT 3.9570 0.8540 4.0070 1.0090 ;
        RECT 3.6230 0.8040 4.0070 0.8540 ;
        RECT 3.6230 0.8540 3.6730 1.5460 ;
        RECT 3.9570 0.3590 4.0070 0.8040 ;
        RECT 3.6230 0.3090 4.0070 0.3590 ;
        RECT 3.6230 0.1480 3.6730 0.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 4.5230 1.7730 ;
    LAYER M1 ;
      RECT 1.1910 0.2990 1.2810 0.3810 ;
      RECT 1.2150 0.3810 1.2650 0.9880 ;
      RECT 0.4310 0.9880 1.2650 1.0380 ;
      RECT 1.1910 1.0380 1.2410 1.3140 ;
      RECT 0.4310 1.0380 0.4810 1.2160 ;
      RECT 0.4310 0.8290 0.4810 0.9880 ;
      RECT 0.4310 0.5790 0.5210 0.6290 ;
      RECT 0.4310 0.4550 0.4810 0.5790 ;
      RECT 0.4310 0.7800 0.5210 0.8290 ;
      RECT 0.4710 0.6290 0.5210 0.7800 ;
      RECT 3.0910 0.0880 3.1410 0.2300 ;
      RECT 2.2490 0.2300 3.1410 0.2800 ;
      RECT 2.4670 0.2800 2.5490 0.3120 ;
      RECT 2.4670 0.2100 2.5490 0.2300 ;
      RECT 2.2490 0.2800 2.2990 0.3140 ;
      RECT 2.0980 0.3140 2.2990 0.3640 ;
      RECT 2.0980 0.3640 2.1480 0.5400 ;
      RECT 1.8590 0.5400 2.1480 0.5900 ;
      RECT 1.3430 0.6400 2.2450 0.6900 ;
      RECT 1.3430 0.6900 1.3930 1.1580 ;
      RECT 1.3430 0.4840 1.3930 0.6400 ;
      RECT 1.3430 1.2080 1.3930 1.3140 ;
      RECT 1.3430 0.3550 1.3930 0.4340 ;
      RECT 1.3430 1.1580 1.7130 1.2080 ;
      RECT 1.3430 0.4340 1.5610 0.4840 ;
      RECT 2.5590 0.4380 3.9010 0.4880 ;
      RECT 3.8510 0.4880 3.9010 0.7040 ;
      RECT 3.5110 0.7040 3.9010 0.7540 ;
      RECT 2.5590 0.4880 2.6090 1.1650 ;
      RECT 2.8620 0.4880 2.9120 0.7660 ;
      RECT 2.8620 0.7660 3.0050 0.8160 ;
      RECT 3.5110 0.7540 3.5610 1.2080 ;
      RECT 3.1510 1.2080 3.5610 1.2580 ;
      RECT 1.8590 0.7860 2.3810 0.8360 ;
      RECT 2.3310 0.6210 2.3810 0.7860 ;
      RECT 2.4070 0.5050 2.4970 0.5550 ;
      RECT 2.4470 0.5550 2.4970 1.0010 ;
      RECT 2.4070 0.4700 2.4570 0.5050 ;
      RECT 1.5500 1.0010 2.4970 1.0510 ;
      RECT 2.2240 0.4200 2.4570 0.4700 ;
      RECT 2.4070 1.0510 2.4570 1.3080 ;
      RECT 2.4070 0.3710 2.4570 0.4200 ;
      RECT 2.2550 1.3080 2.4570 1.3580 ;
      RECT 2.2550 1.1010 2.3050 1.3080 ;
      RECT 1.0850 0.0960 1.4910 0.1460 ;
      RECT 3.0550 0.6040 3.7650 0.6540 ;
      RECT 3.0550 0.6540 3.1050 0.9780 ;
      RECT 2.6940 0.9780 3.1050 1.0280 ;
      RECT 2.6940 0.5880 2.7440 0.9780 ;
      RECT 2.6940 0.5380 2.8010 0.5880 ;
      RECT 1.4190 1.4780 1.9410 1.5280 ;
      RECT 1.4190 1.5280 1.4690 1.5650 ;
      RECT 1.2670 1.4280 1.3170 1.5260 ;
      RECT 1.2670 1.3780 2.0770 1.4280 ;
      RECT 2.0270 1.4280 2.0770 1.5840 ;
      RECT 0.7850 1.5260 1.3170 1.5760 ;
      RECT 0.5830 0.6180 1.0290 0.6680 ;
      RECT 0.5830 0.6680 0.6330 0.9140 ;
      RECT 0.5830 0.4220 0.6330 0.6180 ;
      RECT 1.0390 0.5180 1.1650 0.5680 ;
      RECT 1.0390 0.3940 1.0890 0.5180 ;
      RECT 1.1150 0.5680 1.1650 0.7180 ;
      RECT 1.0390 0.7180 1.1650 0.7680 ;
      RECT 1.0390 0.7680 1.0890 0.9140 ;
      RECT 3.0740 1.4290 3.4610 1.4790 ;
      RECT 3.2380 0.7090 3.4610 0.7590 ;
      RECT 3.2380 0.7590 3.2880 1.0990 ;
      RECT 2.6830 1.0990 3.2880 1.1490 ;
      RECT 2.6830 1.1490 2.7330 1.2720 ;
      RECT 2.5070 1.2720 2.7330 1.3220 ;
      RECT 2.5070 1.3220 2.5570 1.5280 ;
      RECT 2.3150 1.5280 2.5570 1.5780 ;
      RECT 1.4790 1.2780 1.8650 1.3280 ;
    LAYER PO ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 3.7090 0.0680 3.7390 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 4.3170 0.0680 4.3470 1.6060 ;
      RECT 1.2770 0.0680 1.3070 0.5420 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 1.2770 0.7900 1.3070 1.6060 ;
      RECT 3.4050 1.0120 3.4350 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 1.8850 0.0680 1.9150 0.6180 ;
      RECT 3.4050 0.0680 3.4350 0.7870 ;
      RECT 2.4930 0.8250 2.5230 1.6060 ;
      RECT 2.4930 0.0680 2.5230 0.6220 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 1.8850 0.7580 1.9150 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
  END
END DFFNARX1_LVT

MACRO DFFNARX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.56 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.7750 0.8040 4.3210 0.8540 ;
        RECT 3.7750 0.8540 3.8250 1.5460 ;
        RECT 4.2710 0.5110 4.3210 0.8040 ;
        RECT 4.2010 0.4510 4.3210 0.5110 ;
        RECT 3.7750 0.4010 4.3210 0.4510 ;
        RECT 3.7750 0.1480 3.8250 0.4010 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.3530 0.2490 4.4630 0.2700 ;
        RECT 4.0790 0.2700 4.4630 0.3200 ;
        RECT 4.3530 0.3200 4.4630 0.3590 ;
        RECT 4.0790 0.1480 4.1290 0.2700 ;
        RECT 4.3950 0.3590 4.4450 0.9180 ;
        RECT 4.0790 0.9180 4.4450 0.9680 ;
        RECT 4.0790 0.9680 4.1290 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.5600 0.0300 ;
        RECT 0.5860 0.0300 0.6360 0.1960 ;
        RECT 4.2310 0.0300 4.2810 0.2200 ;
        RECT 3.9270 0.0300 3.9770 0.3190 ;
        RECT 3.6230 0.0300 3.6730 0.4080 ;
        RECT 0.2790 0.0300 0.3290 0.4190 ;
        RECT 1.5410 0.0300 1.5910 0.2870 ;
        RECT 3.4710 0.0300 3.5210 0.3300 ;
        RECT 0.5860 0.1960 0.9370 0.2460 ;
        RECT 1.5410 0.2870 2.0010 0.3370 ;
        RECT 2.9990 0.3300 3.5370 0.3800 ;
        RECT 0.8870 0.2460 0.9370 0.4500 ;
        RECT 0.7350 0.2460 0.7850 0.4500 ;
        RECT 1.9510 0.3370 2.0010 0.4610 ;
        RECT 1.9510 0.2490 2.0010 0.2870 ;
        RECT 1.9510 0.1990 2.1760 0.2490 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.5600 1.7020 ;
        RECT 0.2790 1.0330 0.3290 1.6420 ;
        RECT 3.6230 0.9120 3.6730 1.6420 ;
        RECT 4.2310 1.0520 4.2810 1.6420 ;
        RECT 3.9270 0.9600 3.9770 1.6420 ;
        RECT 3.5110 1.3580 3.5610 1.6420 ;
        RECT 2.1270 1.3280 2.1770 1.6420 ;
        RECT 0.4330 1.3640 0.4830 1.6420 ;
        RECT 2.8340 1.3080 3.5610 1.3580 ;
        RECT 1.9340 1.2780 2.1770 1.3280 ;
        RECT 0.4330 1.3440 0.9370 1.3640 ;
        RECT 0.4340 1.3140 0.9370 1.3440 ;
        RECT 0.7350 1.0980 0.7850 1.3140 ;
        RECT 0.8870 1.1110 0.9370 1.3140 ;
    END
  END VDD

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7230 0.0900 2.8530 0.1400 ;
        RECT 2.7710 0.1400 2.8530 0.1760 ;
        RECT 1.7230 0.1400 1.8790 0.2190 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.3590 0.6800 ;
        RECT 0.2490 0.6800 0.4210 0.7300 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.4240 0.7250 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 4.6760 1.7730 ;
    LAYER M1 ;
      RECT 1.1910 0.2990 1.2810 0.3810 ;
      RECT 1.2150 0.3810 1.2650 0.9880 ;
      RECT 0.4310 0.9880 1.2650 1.0380 ;
      RECT 1.1910 1.0380 1.2410 1.3140 ;
      RECT 0.4310 1.0380 0.4810 1.2160 ;
      RECT 0.4310 0.8290 0.4810 0.9880 ;
      RECT 0.4310 0.5790 0.5210 0.6290 ;
      RECT 0.4310 0.4550 0.4810 0.5790 ;
      RECT 0.4310 0.7800 0.5210 0.8290 ;
      RECT 0.4710 0.6290 0.5210 0.7800 ;
      RECT 3.0910 0.1020 3.1410 0.2300 ;
      RECT 2.2490 0.2300 3.1410 0.2800 ;
      RECT 2.4670 0.1980 2.5490 0.2300 ;
      RECT 2.2490 0.2800 2.2990 0.3140 ;
      RECT 2.0980 0.3140 2.2990 0.3640 ;
      RECT 2.0980 0.3640 2.1480 0.5860 ;
      RECT 1.8590 0.5860 2.1480 0.6360 ;
      RECT 1.3430 0.6860 2.2450 0.7360 ;
      RECT 1.3430 0.7360 1.3930 1.1580 ;
      RECT 1.3430 0.4840 1.3930 0.6860 ;
      RECT 1.3430 1.2080 1.3930 1.3140 ;
      RECT 1.3430 0.3550 1.3930 0.4340 ;
      RECT 1.3430 1.1580 1.7130 1.2080 ;
      RECT 1.3430 0.4340 1.5610 0.4840 ;
      RECT 3.9840 0.6040 4.2210 0.6540 ;
      RECT 2.8620 0.4880 2.9120 0.5030 ;
      RECT 2.8620 0.5530 2.9120 0.7660 ;
      RECT 3.5110 0.7540 3.5610 1.2080 ;
      RECT 2.5590 0.4380 2.9120 0.4880 ;
      RECT 2.8620 0.7660 3.0050 0.8160 ;
      RECT 3.1510 1.2080 3.5610 1.2580 ;
      RECT 2.5590 0.4880 2.6090 1.1650 ;
      RECT 3.9840 0.5530 4.0340 0.6040 ;
      RECT 3.9840 0.6540 4.0340 0.7040 ;
      RECT 2.8620 0.5030 4.0340 0.5530 ;
      RECT 3.5110 0.7040 4.0340 0.7540 ;
      RECT 1.8590 0.7860 2.3810 0.8360 ;
      RECT 2.3310 0.6210 2.3810 0.7860 ;
      RECT 2.4070 0.5050 2.4970 0.5550 ;
      RECT 2.4470 0.5550 2.4970 1.0010 ;
      RECT 2.4070 0.4700 2.4570 0.5050 ;
      RECT 1.5500 1.0010 2.4970 1.0510 ;
      RECT 2.2240 0.4200 2.4570 0.4700 ;
      RECT 2.4070 1.0510 2.4570 1.3080 ;
      RECT 2.4070 0.3710 2.4570 0.4200 ;
      RECT 2.2550 1.3080 2.4570 1.3580 ;
      RECT 2.2550 1.1010 2.3050 1.3080 ;
      RECT 1.0850 0.0960 1.4910 0.1460 ;
      RECT 3.0550 0.6040 3.9170 0.6540 ;
      RECT 3.0550 0.6540 3.1050 0.9780 ;
      RECT 2.6940 0.9780 3.1050 1.0280 ;
      RECT 2.6940 0.5880 2.7440 0.9780 ;
      RECT 2.6940 0.5380 2.8010 0.5880 ;
      RECT 1.4190 1.4780 1.9410 1.5280 ;
      RECT 1.4190 1.5280 1.4690 1.5650 ;
      RECT 1.2670 1.4280 1.3170 1.5260 ;
      RECT 1.2670 1.3780 2.0770 1.4280 ;
      RECT 2.0270 1.4280 2.0770 1.5740 ;
      RECT 0.7850 1.5260 1.3170 1.5760 ;
      RECT 0.5830 0.6180 1.0290 0.6680 ;
      RECT 0.5830 0.6680 0.6330 0.9140 ;
      RECT 0.5830 0.4220 0.6330 0.6180 ;
      RECT 1.0390 0.5180 1.1650 0.5680 ;
      RECT 1.0390 0.3940 1.0890 0.5180 ;
      RECT 1.1150 0.5680 1.1650 0.7180 ;
      RECT 1.0390 0.7180 1.1650 0.7680 ;
      RECT 1.0390 0.7680 1.0890 0.9140 ;
      RECT 3.0740 1.4290 3.4610 1.4790 ;
      RECT 3.2380 0.7090 3.4610 0.7590 ;
      RECT 3.2380 0.7590 3.2880 1.0990 ;
      RECT 2.6830 1.0990 3.2880 1.1490 ;
      RECT 2.6830 1.1490 2.7330 1.2720 ;
      RECT 2.5070 1.2720 2.7330 1.3220 ;
      RECT 2.5070 1.3220 2.5570 1.5280 ;
      RECT 2.3150 1.5280 2.5570 1.5780 ;
      RECT 1.4790 1.2780 1.8650 1.3280 ;
    LAYER PO ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 1.8850 0.7580 1.9150 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 1.2770 0.0680 1.3070 0.5420 ;
      RECT 1.2770 0.7900 1.3070 1.6060 ;
      RECT 3.4050 1.0120 3.4350 1.6060 ;
      RECT 4.3170 0.0680 4.3470 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 4.4690 0.0680 4.4990 1.6060 ;
      RECT 1.8850 0.0680 1.9150 0.6410 ;
      RECT 3.4050 0.0680 3.4350 0.7870 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 2.4930 0.8250 2.5230 1.6060 ;
      RECT 3.7090 0.0680 3.7390 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 2.4930 0.0680 2.5230 0.6220 ;
  END
END DFFNARX2_LVT

MACRO DFFNASRNX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.408 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.4080 0.0300 ;
        RECT 0.5860 0.0300 0.6360 0.1960 ;
        RECT 0.2790 0.0300 0.3290 0.4190 ;
        RECT 3.9270 0.0300 3.9770 0.2200 ;
        RECT 3.7750 0.0300 3.8250 0.3300 ;
        RECT 1.5410 0.0300 1.5910 0.2870 ;
        RECT 0.5860 0.1960 0.9370 0.2460 ;
        RECT 3.1510 0.3300 3.8410 0.3800 ;
        RECT 1.5410 0.2870 2.1530 0.3370 ;
        RECT 0.8870 0.2460 0.9370 0.4500 ;
        RECT 0.7350 0.2460 0.7850 0.4500 ;
        RECT 2.1030 0.3370 2.1530 0.4610 ;
        RECT 1.9510 0.3370 2.0010 0.4610 ;
    END
  END VSS

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0490 0.8570 4.1600 0.9670 ;
        RECT 4.1030 0.2040 4.1530 0.8570 ;
        RECT 4.1030 0.9670 4.1530 1.2210 ;
        RECT 4.0630 0.1540 4.1530 0.2040 ;
        RECT 4.0790 1.2210 4.1530 1.2710 ;
        RECT 4.0790 1.2710 4.1290 1.5460 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.4080 1.7020 ;
        RECT 0.2790 1.0330 0.3290 1.6420 ;
        RECT 3.9270 0.9470 3.9770 1.6420 ;
        RECT 2.1270 1.3280 2.1770 1.6420 ;
        RECT 3.8150 1.3580 3.8650 1.6420 ;
        RECT 0.4330 1.3580 0.4830 1.6420 ;
        RECT 1.9340 1.2780 2.3360 1.3280 ;
        RECT 2.9860 1.3080 3.8650 1.3580 ;
        RECT 0.4330 1.3380 0.9370 1.3580 ;
        RECT 0.4340 1.3080 0.9370 1.3380 ;
        RECT 0.7350 1.0920 0.7850 1.3080 ;
        RECT 0.8870 1.1050 0.9370 1.3080 ;
    END
  END VDD

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7230 0.0880 3.0050 0.1380 ;
        RECT 2.9230 0.1380 3.0050 0.1740 ;
        RECT 1.7230 0.1380 1.8790 0.2070 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.3590 0.6800 ;
        RECT 0.2490 0.6800 0.4210 0.7300 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.5310 0.8570 3.7030 1.0340 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.4240 0.7250 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 4.5230 1.7730 ;
    LAYER M1 ;
      RECT 1.8590 0.8820 2.5330 0.9320 ;
      RECT 2.4830 0.5970 2.5330 0.8820 ;
      RECT 1.1910 0.2990 1.2810 0.3810 ;
      RECT 1.2150 0.3810 1.2650 0.9880 ;
      RECT 0.4310 0.9880 1.2650 1.0380 ;
      RECT 1.1910 1.0380 1.2410 1.3140 ;
      RECT 0.4310 1.0380 0.4810 1.2160 ;
      RECT 0.4310 0.8290 0.4810 0.9880 ;
      RECT 0.4310 0.5790 0.5210 0.6290 ;
      RECT 0.4310 0.4550 0.4810 0.5790 ;
      RECT 0.4310 0.7800 0.5210 0.8290 ;
      RECT 0.4710 0.6290 0.5210 0.7800 ;
      RECT 3.2430 0.0880 3.2930 0.2300 ;
      RECT 2.2950 0.2300 3.2930 0.2800 ;
      RECT 2.6190 0.2800 2.7010 0.3010 ;
      RECT 2.6190 0.1990 2.7010 0.2300 ;
      RECT 2.2950 0.2800 2.3450 0.5840 ;
      RECT 1.8590 0.5840 2.3450 0.6340 ;
      RECT 1.3430 0.6840 2.2450 0.7340 ;
      RECT 1.3430 0.7340 1.3930 1.1580 ;
      RECT 1.3430 0.4840 1.3930 0.6840 ;
      RECT 1.3430 1.2080 1.3930 1.3140 ;
      RECT 1.3430 0.3550 1.3930 0.4340 ;
      RECT 1.3430 1.1580 1.7130 1.2080 ;
      RECT 1.3430 0.4340 1.5610 0.4840 ;
      RECT 3.8150 0.7040 4.0530 0.7540 ;
      RECT 4.0030 0.4880 4.0530 0.7040 ;
      RECT 2.7110 0.4380 4.0530 0.4880 ;
      RECT 3.8150 0.7540 3.8650 1.1080 ;
      RECT 3.4550 1.1080 3.8650 1.1580 ;
      RECT 2.7110 0.4880 2.7610 1.1650 ;
      RECT 3.0140 0.4880 3.0640 0.7660 ;
      RECT 3.0140 0.7660 3.1570 0.8160 ;
      RECT 3.2070 0.6040 3.4610 0.6540 ;
      RECT 3.2070 0.6540 3.2570 0.9780 ;
      RECT 2.8460 0.9780 3.2570 1.0280 ;
      RECT 2.8460 0.5880 2.8960 0.9780 ;
      RECT 2.8460 0.5380 2.9530 0.5880 ;
      RECT 1.5500 1.0010 2.6490 1.0510 ;
      RECT 2.5990 0.4960 2.6490 1.0010 ;
      RECT 2.5590 1.0510 2.6090 1.3080 ;
      RECT 2.4070 0.4460 2.6490 0.4960 ;
      RECT 2.4070 1.3080 2.6090 1.3580 ;
      RECT 2.5590 0.3710 2.6090 0.4460 ;
      RECT 2.4070 0.3710 2.4570 0.4460 ;
      RECT 2.4070 1.2160 2.4570 1.3080 ;
      RECT 2.0860 1.1660 2.4570 1.2160 ;
      RECT 3.2260 1.4080 3.7650 1.4580 ;
      RECT 1.4190 1.4780 1.9410 1.5280 ;
      RECT 1.4190 1.5280 1.4690 1.5650 ;
      RECT 0.7950 1.5260 1.3170 1.5760 ;
      RECT 1.2670 1.4280 1.3170 1.5260 ;
      RECT 1.2670 1.3780 2.0770 1.4280 ;
      RECT 2.0270 1.4280 2.0770 1.5440 ;
      RECT 0.5830 0.6180 1.0290 0.6680 ;
      RECT 0.5830 0.6680 0.6330 0.9140 ;
      RECT 0.5830 0.4220 0.6330 0.6180 ;
      RECT 1.0390 0.5180 1.1650 0.5680 ;
      RECT 1.0390 0.3940 1.0890 0.5180 ;
      RECT 1.1150 0.5680 1.1650 0.7180 ;
      RECT 1.0390 0.7180 1.1650 0.7680 ;
      RECT 1.0390 0.7680 1.0890 0.9140 ;
      RECT 3.3450 0.7090 3.7650 0.7590 ;
      RECT 3.3450 0.7590 3.3950 1.0990 ;
      RECT 2.8350 1.0990 3.3950 1.1490 ;
      RECT 2.8350 1.1490 2.8850 1.2720 ;
      RECT 2.6590 1.2720 2.8850 1.3220 ;
      RECT 2.6590 1.3220 2.7090 1.4280 ;
      RECT 2.4670 1.4280 2.7090 1.4780 ;
      RECT 1.0990 0.0960 1.4910 0.1460 ;
      RECT 2.2860 1.5280 3.6260 1.5780 ;
      RECT 3.3030 1.2080 3.6890 1.2580 ;
      RECT 1.4790 1.2780 1.8650 1.3280 ;
    LAYER PO ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 1.2770 0.0680 1.3070 0.5420 ;
      RECT 1.2770 0.7900 1.3070 1.6060 ;
      RECT 3.7090 0.0680 3.7390 0.7870 ;
      RECT 1.8850 0.0680 1.9150 0.6620 ;
      RECT 3.7090 1.0120 3.7390 1.6060 ;
      RECT 2.6450 0.7320 2.6750 1.6060 ;
      RECT 2.6450 0.0680 2.6750 0.6220 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 1.8850 0.8540 1.9150 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 4.3170 0.0680 4.3470 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
  END
END DFFNASRNX1_LVT

MACRO DFFNASRNX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.56 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.5600 0.0300 ;
        RECT 0.5860 0.0300 0.6360 0.1960 ;
        RECT 3.9270 0.0300 3.9770 0.5060 ;
        RECT 4.2310 0.0300 4.2810 0.3120 ;
        RECT 0.2790 0.0300 0.3290 0.4190 ;
        RECT 3.7750 0.0300 3.8250 0.3300 ;
        RECT 1.5410 0.0300 1.5910 0.2870 ;
        RECT 0.5860 0.1960 0.9370 0.2460 ;
        RECT 3.1510 0.3300 3.8410 0.3800 ;
        RECT 1.5410 0.2870 2.1530 0.3370 ;
        RECT 0.8870 0.2460 0.9370 0.4500 ;
        RECT 0.7350 0.2460 0.7850 0.4500 ;
        RECT 2.1030 0.3370 2.1530 0.4610 ;
        RECT 1.9510 0.3370 2.0010 0.4610 ;
    END
  END VSS

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0790 0.7650 4.4630 0.8150 ;
        RECT 4.0790 0.8150 4.1290 1.5460 ;
        RECT 4.3090 0.7050 4.4630 0.7650 ;
        RECT 4.3090 0.5130 4.3590 0.7050 ;
        RECT 4.0790 0.4630 4.3590 0.5130 ;
        RECT 4.0790 0.1380 4.1290 0.4630 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.5600 1.7020 ;
        RECT 0.2790 1.0330 0.3290 1.6420 ;
        RECT 3.9270 0.9220 3.9770 1.6420 ;
        RECT 4.2310 0.9220 4.2810 1.6420 ;
        RECT 2.1270 1.3280 2.1770 1.6420 ;
        RECT 3.8150 1.3580 3.8650 1.6420 ;
        RECT 0.4330 1.3580 0.4830 1.6420 ;
        RECT 1.9340 1.2780 2.3360 1.3280 ;
        RECT 2.9860 1.3080 3.8650 1.3580 ;
        RECT 0.4330 1.3380 0.9370 1.3580 ;
        RECT 0.4340 1.3080 0.9370 1.3380 ;
        RECT 0.7350 1.0920 0.7850 1.3080 ;
        RECT 0.8870 1.1050 0.9370 1.3080 ;
    END
  END VDD

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9230 0.1380 3.0050 0.1740 ;
        RECT 1.7230 0.0880 3.0050 0.1380 ;
        RECT 1.7230 0.1380 1.8790 0.2070 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.3590 0.6800 ;
        RECT 0.2490 0.6800 0.4210 0.7300 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.5310 0.8570 3.7030 1.0340 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.4240 0.7250 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 4.6750 1.7730 ;
    LAYER M1 ;
      RECT 1.8590 0.8820 2.5330 0.9320 ;
      RECT 2.4830 0.5970 2.5330 0.8820 ;
      RECT 1.1910 0.2990 1.2810 0.3810 ;
      RECT 1.2150 0.3810 1.2650 0.9880 ;
      RECT 0.4310 0.9880 1.2650 1.0380 ;
      RECT 1.1910 1.0380 1.2410 1.3140 ;
      RECT 0.4310 1.0380 0.4810 1.2160 ;
      RECT 0.4310 0.8290 0.4810 0.9880 ;
      RECT 0.4310 0.5790 0.5210 0.6290 ;
      RECT 0.4310 0.4550 0.4810 0.5790 ;
      RECT 0.4310 0.7800 0.5210 0.8290 ;
      RECT 0.4710 0.6290 0.5210 0.7800 ;
      RECT 3.2430 0.0880 3.2930 0.2300 ;
      RECT 2.2950 0.2300 3.2930 0.2800 ;
      RECT 2.6190 0.2800 2.7010 0.2900 ;
      RECT 2.2950 0.2800 2.3450 0.5840 ;
      RECT 1.8590 0.5840 2.3450 0.6340 ;
      RECT 2.6190 0.1880 2.7010 0.2300 ;
      RECT 1.3430 0.6840 2.2450 0.7340 ;
      RECT 1.3430 0.7340 1.3930 1.1580 ;
      RECT 1.3430 0.4840 1.3930 0.6840 ;
      RECT 1.3430 1.2080 1.3930 1.3140 ;
      RECT 1.3430 0.3550 1.3930 0.4340 ;
      RECT 1.3430 1.1580 1.7130 1.2080 ;
      RECT 1.3430 0.4340 1.5610 0.4840 ;
      RECT 3.8150 0.6040 4.2210 0.6540 ;
      RECT 3.8150 0.6540 3.8650 1.1080 ;
      RECT 3.8150 0.4880 3.8650 0.6040 ;
      RECT 3.4550 1.1080 3.8650 1.1580 ;
      RECT 2.7110 0.4380 3.8650 0.4880 ;
      RECT 2.7110 0.4880 2.7610 1.1650 ;
      RECT 3.0140 0.4880 3.0640 0.7660 ;
      RECT 3.0140 0.7660 3.1570 0.8160 ;
      RECT 1.5500 1.0010 2.6490 1.0510 ;
      RECT 2.5990 0.4960 2.6490 1.0010 ;
      RECT 2.5590 1.0510 2.6090 1.3080 ;
      RECT 2.4070 0.4460 2.6490 0.4960 ;
      RECT 2.4070 1.3080 2.6090 1.3580 ;
      RECT 2.5590 0.3710 2.6090 0.4460 ;
      RECT 2.4070 0.3710 2.4570 0.4460 ;
      RECT 2.4070 1.2160 2.4570 1.3080 ;
      RECT 2.0860 1.1660 2.4570 1.2160 ;
      RECT 3.2070 0.6040 3.4610 0.6540 ;
      RECT 3.2070 0.6540 3.2570 0.9780 ;
      RECT 2.8460 0.9780 3.2570 1.0280 ;
      RECT 2.8460 0.5880 2.8960 0.9780 ;
      RECT 2.8460 0.5380 2.9530 0.5880 ;
      RECT 3.2260 1.4080 3.7650 1.4580 ;
      RECT 1.4190 1.4780 1.9410 1.5280 ;
      RECT 1.4190 1.5280 1.4690 1.5650 ;
      RECT 0.7950 1.5260 1.3170 1.5760 ;
      RECT 1.2670 1.4280 1.3170 1.5260 ;
      RECT 1.2670 1.3780 2.0770 1.4280 ;
      RECT 2.0270 1.4280 2.0770 1.5440 ;
      RECT 0.5830 0.6180 1.0290 0.6680 ;
      RECT 0.5830 0.6680 0.6330 0.9140 ;
      RECT 0.5830 0.4220 0.6330 0.6180 ;
      RECT 1.0390 0.5180 1.1650 0.5680 ;
      RECT 1.0390 0.3940 1.0890 0.5180 ;
      RECT 1.1150 0.5680 1.1650 0.7180 ;
      RECT 1.0390 0.7180 1.1650 0.7680 ;
      RECT 1.0390 0.7680 1.0890 0.9140 ;
      RECT 3.3450 0.7090 3.7650 0.7590 ;
      RECT 3.3450 0.7590 3.3950 1.0990 ;
      RECT 2.8350 1.0990 3.3950 1.1490 ;
      RECT 2.8350 1.1490 2.8850 1.2720 ;
      RECT 2.6590 1.2720 2.8850 1.3220 ;
      RECT 2.6590 1.3220 2.7090 1.4280 ;
      RECT 2.4670 1.4280 2.7090 1.4780 ;
      RECT 1.0990 0.0960 1.4910 0.1460 ;
      RECT 2.2860 1.5280 3.6260 1.5780 ;
      RECT 3.3030 1.2080 3.6890 1.2580 ;
      RECT 1.4790 1.2780 1.8650 1.3280 ;
    LAYER PO ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 1.2770 0.0680 1.3070 0.5420 ;
      RECT 1.2770 0.7900 1.3070 1.6060 ;
      RECT 3.7090 0.0680 3.7390 0.7870 ;
      RECT 1.8850 0.0680 1.9150 0.6620 ;
      RECT 4.4690 0.0680 4.4990 1.6060 ;
      RECT 3.7090 1.0120 3.7390 1.6060 ;
      RECT 2.6450 0.7320 2.6750 1.6060 ;
      RECT 2.6450 0.0680 2.6750 0.6220 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 1.8850 0.8540 1.9150 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 4.3170 0.0680 4.3470 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
  END
END DFFNASRNX2_LVT

MACRO DFFNASRQX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.408 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.4080 0.0300 ;
        RECT 0.5860 0.0300 0.6360 0.1960 ;
        RECT 0.2790 0.0300 0.3290 0.4190 ;
        RECT 4.0790 0.0300 4.1290 0.2200 ;
        RECT 3.7750 0.0300 3.8250 0.3300 ;
        RECT 1.5410 0.0300 1.5910 0.2870 ;
        RECT 0.5860 0.1960 0.9370 0.2460 ;
        RECT 3.1510 0.3300 3.8410 0.3800 ;
        RECT 1.5410 0.2870 2.1530 0.3370 ;
        RECT 0.8870 0.2460 0.9370 0.4500 ;
        RECT 0.7350 0.2460 0.7850 0.4500 ;
        RECT 2.1030 0.3370 2.1530 0.4610 ;
        RECT 1.9510 0.3370 2.0010 0.4610 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.4080 1.7020 ;
        RECT 0.2790 1.0330 0.3290 1.6420 ;
        RECT 4.0790 0.9470 4.1290 1.6420 ;
        RECT 2.1270 1.3280 2.1770 1.6420 ;
        RECT 3.8150 1.3580 3.8650 1.6420 ;
        RECT 0.4330 1.3580 0.4830 1.6420 ;
        RECT 1.9340 1.2780 2.3360 1.3280 ;
        RECT 2.9860 1.3080 3.8650 1.3580 ;
        RECT 0.4330 1.3380 0.9370 1.3580 ;
        RECT 0.4340 1.3080 0.9370 1.3380 ;
        RECT 0.7350 1.0920 0.7850 1.3080 ;
        RECT 0.8870 1.1050 0.9370 1.3080 ;
    END
  END VDD

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9230 0.1380 3.0050 0.1740 ;
        RECT 1.7230 0.0880 3.0050 0.1380 ;
        RECT 1.7230 0.1380 1.8790 0.2070 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.3590 0.6800 ;
        RECT 0.2490 0.6800 0.4210 0.7300 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.5310 0.8570 3.7030 1.0340 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.4240 0.7250 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.2010 1.0090 4.3110 1.1190 ;
        RECT 4.2190 0.8540 4.2690 1.0090 ;
        RECT 3.9270 0.8040 4.2690 0.8540 ;
        RECT 3.9270 0.8540 3.9770 1.5460 ;
        RECT 4.2190 0.3590 4.2690 0.8040 ;
        RECT 3.9270 0.3090 4.2690 0.3590 ;
        RECT 3.9270 0.1480 3.9770 0.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 4.5230 1.7730 ;
    LAYER M1 ;
      RECT 1.1910 0.2990 1.2810 0.3810 ;
      RECT 1.2150 0.3810 1.2650 0.9880 ;
      RECT 0.4310 0.9880 1.2650 1.0380 ;
      RECT 1.1910 1.0380 1.2410 1.3140 ;
      RECT 0.4310 1.0380 0.4810 1.2160 ;
      RECT 0.4310 0.8290 0.4810 0.9880 ;
      RECT 0.4310 0.5790 0.5210 0.6290 ;
      RECT 0.4310 0.4550 0.4810 0.5790 ;
      RECT 0.4310 0.7800 0.5210 0.8290 ;
      RECT 0.4710 0.6290 0.5210 0.7800 ;
      RECT 3.2430 0.0880 3.2930 0.2300 ;
      RECT 2.2950 0.2300 3.2930 0.2800 ;
      RECT 2.6190 0.2800 2.7010 0.3020 ;
      RECT 2.6190 0.2000 2.7010 0.2300 ;
      RECT 2.2950 0.2800 2.3450 0.5890 ;
      RECT 1.8590 0.5890 2.3450 0.6390 ;
      RECT 1.3430 0.6890 2.2450 0.7390 ;
      RECT 1.3430 0.4840 1.3930 0.6890 ;
      RECT 1.3430 0.7390 1.3930 1.1580 ;
      RECT 1.3430 0.3550 1.3930 0.4340 ;
      RECT 1.3430 1.2080 1.3930 1.3140 ;
      RECT 1.3430 0.4340 1.5610 0.4840 ;
      RECT 1.3430 1.1580 1.7130 1.2080 ;
      RECT 4.1190 0.4880 4.1690 0.7040 ;
      RECT 2.7110 0.4380 4.1690 0.4880 ;
      RECT 3.8150 0.7040 4.1690 0.7540 ;
      RECT 3.8150 0.7540 3.8650 1.1080 ;
      RECT 3.4550 1.1080 3.8650 1.1580 ;
      RECT 2.7110 0.4880 2.7610 1.1650 ;
      RECT 3.0140 0.4880 3.0640 0.7660 ;
      RECT 3.0140 0.7660 3.1570 0.8160 ;
      RECT 1.8590 0.8870 2.5330 0.9370 ;
      RECT 2.4830 0.6020 2.5330 0.8870 ;
      RECT 1.5500 1.0010 2.6490 1.0510 ;
      RECT 2.5990 0.4960 2.6490 1.0010 ;
      RECT 2.5590 1.0510 2.6090 1.3080 ;
      RECT 2.4070 0.4460 2.6490 0.4960 ;
      RECT 2.4070 1.3080 2.6090 1.3580 ;
      RECT 2.5590 0.3710 2.6090 0.4460 ;
      RECT 2.4070 0.3710 2.4570 0.4460 ;
      RECT 2.4070 1.2160 2.4570 1.3080 ;
      RECT 2.0860 1.1660 2.4570 1.2160 ;
      RECT 3.2070 0.6040 4.0690 0.6540 ;
      RECT 3.2070 0.6540 3.2570 0.9780 ;
      RECT 2.8460 0.9780 3.2570 1.0280 ;
      RECT 2.8460 0.5880 2.8960 0.9780 ;
      RECT 2.8460 0.5380 2.9530 0.5880 ;
      RECT 3.2260 1.4080 3.7650 1.4580 ;
      RECT 1.4190 1.4780 1.9410 1.5280 ;
      RECT 1.4190 1.5280 1.4690 1.5650 ;
      RECT 0.7950 1.5260 1.3170 1.5760 ;
      RECT 1.2670 1.4280 1.3170 1.5260 ;
      RECT 1.2670 1.3780 2.0770 1.4280 ;
      RECT 2.0270 1.4280 2.0770 1.5440 ;
      RECT 0.5830 0.6180 1.0290 0.6680 ;
      RECT 0.5830 0.6680 0.6330 0.9140 ;
      RECT 0.5830 0.4220 0.6330 0.6180 ;
      RECT 1.0390 0.5180 1.1650 0.5680 ;
      RECT 1.0390 0.3940 1.0890 0.5180 ;
      RECT 1.1150 0.5680 1.1650 0.7180 ;
      RECT 1.0390 0.7180 1.1650 0.7680 ;
      RECT 1.0390 0.7680 1.0890 0.9140 ;
      RECT 3.3450 0.7090 3.7650 0.7590 ;
      RECT 3.3450 0.7590 3.3950 1.0990 ;
      RECT 2.8350 1.0990 3.3950 1.1490 ;
      RECT 2.8350 1.1490 2.8850 1.2720 ;
      RECT 2.6590 1.2720 2.8850 1.3220 ;
      RECT 2.6590 1.3220 2.7090 1.4280 ;
      RECT 2.4670 1.4280 2.7090 1.4780 ;
      RECT 1.0990 0.0960 1.4910 0.1460 ;
      RECT 2.2860 1.5280 3.6260 1.5780 ;
      RECT 3.3030 1.2080 3.6890 1.2580 ;
      RECT 1.4790 1.2780 1.8650 1.3280 ;
    LAYER PO ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 1.2770 0.0680 1.3070 0.5420 ;
      RECT 3.7090 0.0680 3.7390 0.7870 ;
      RECT 2.6450 0.0680 2.6750 0.6220 ;
      RECT 1.8850 0.8530 1.9150 1.6060 ;
      RECT 1.8850 0.0680 1.9150 0.6610 ;
      RECT 2.6450 0.7320 2.6750 1.6060 ;
      RECT 3.7090 1.0120 3.7390 1.6060 ;
      RECT 1.2770 0.7900 1.3070 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 4.3170 0.0680 4.3470 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
  END
END DFFNASRQX1_LVT

MACRO DFFNASRQX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.56 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.5600 0.0300 ;
        RECT 0.5860 0.0300 0.6360 0.1960 ;
        RECT 0.2790 0.0300 0.3290 0.4190 ;
        RECT 3.9270 0.0300 3.9770 0.4150 ;
        RECT 4.2310 0.0300 4.2810 0.3120 ;
        RECT 3.7750 0.0300 3.8250 0.3300 ;
        RECT 1.5410 0.0300 1.5910 0.2870 ;
        RECT 0.5860 0.1960 0.9370 0.2460 ;
        RECT 3.1510 0.3300 3.8410 0.3800 ;
        RECT 1.5410 0.2870 2.1530 0.3370 ;
        RECT 0.8870 0.2460 0.9370 0.4500 ;
        RECT 0.7350 0.2460 0.7850 0.4500 ;
        RECT 2.1030 0.3370 2.1530 0.4610 ;
        RECT 1.9510 0.3370 2.0010 0.4610 ;
    END
  END VSS

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.3520 0.2490 4.4630 0.3620 ;
        RECT 4.0790 0.3620 4.4210 0.4120 ;
        RECT 4.0790 0.1380 4.1290 0.3620 ;
        RECT 4.3710 0.4120 4.4210 0.8130 ;
        RECT 4.0790 0.8130 4.4210 0.8630 ;
        RECT 4.0790 0.8630 4.1290 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.5600 1.7020 ;
        RECT 0.2790 1.0330 0.3290 1.6420 ;
        RECT 3.9270 0.9220 3.9770 1.6420 ;
        RECT 4.2310 0.9220 4.2810 1.6420 ;
        RECT 2.1270 1.3280 2.1770 1.6420 ;
        RECT 3.8150 1.3580 3.8650 1.6420 ;
        RECT 0.4330 1.3580 0.4830 1.6420 ;
        RECT 1.9340 1.2780 2.3360 1.3280 ;
        RECT 2.9860 1.3080 3.8650 1.3580 ;
        RECT 0.4330 1.3380 0.9370 1.3580 ;
        RECT 0.4340 1.3080 0.9370 1.3380 ;
        RECT 0.7350 1.0920 0.7850 1.3080 ;
        RECT 0.8870 1.1050 0.9370 1.3080 ;
    END
  END VDD

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9230 0.1380 3.0050 0.1740 ;
        RECT 1.7230 0.0880 3.0050 0.1380 ;
        RECT 1.7230 0.1380 1.8790 0.2070 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.3590 0.6800 ;
        RECT 0.2490 0.6800 0.4210 0.7300 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.5310 0.8570 3.7030 1.0340 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.4240 0.7250 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 4.6750 1.7730 ;
    LAYER M1 ;
      RECT 1.1910 0.2990 1.2810 0.3810 ;
      RECT 1.2150 0.3810 1.2650 0.9880 ;
      RECT 0.4310 0.9880 1.2650 1.0380 ;
      RECT 1.1910 1.0380 1.2410 1.3140 ;
      RECT 0.4310 1.0380 0.4810 1.2160 ;
      RECT 0.4310 0.8290 0.4810 0.9880 ;
      RECT 0.4310 0.5790 0.5210 0.6290 ;
      RECT 0.4310 0.4550 0.4810 0.5790 ;
      RECT 0.4310 0.7800 0.5210 0.8290 ;
      RECT 0.4710 0.6290 0.5210 0.7800 ;
      RECT 3.2430 0.0880 3.2930 0.2300 ;
      RECT 2.2950 0.2300 3.2930 0.2800 ;
      RECT 2.6190 0.2800 2.7010 0.2900 ;
      RECT 2.2950 0.2800 2.3450 0.5890 ;
      RECT 1.8590 0.5890 2.3450 0.6390 ;
      RECT 2.6190 0.1880 2.7010 0.2300 ;
      RECT 1.3430 0.6890 2.2450 0.7390 ;
      RECT 1.3430 0.4840 1.3930 0.6890 ;
      RECT 1.3430 0.7390 1.3930 1.1580 ;
      RECT 1.3430 0.3550 1.3930 0.4340 ;
      RECT 1.3430 1.2080 1.3930 1.3140 ;
      RECT 1.3430 0.4340 1.5610 0.4840 ;
      RECT 1.3430 1.1580 1.7130 1.2080 ;
      RECT 3.0140 0.4940 4.3210 0.5440 ;
      RECT 4.2710 0.5440 4.3210 0.7040 ;
      RECT 3.8150 0.7040 4.3210 0.7540 ;
      RECT 3.8150 0.7540 3.8650 1.1080 ;
      RECT 3.4550 1.1080 3.8650 1.1580 ;
      RECT 3.0140 0.5440 3.0640 0.7660 ;
      RECT 3.0140 0.4880 3.0640 0.4940 ;
      RECT 3.0140 0.7660 3.1570 0.8160 ;
      RECT 2.7110 0.4380 3.0640 0.4880 ;
      RECT 2.7110 0.4880 2.7610 1.1650 ;
      RECT 1.8590 0.8870 2.5330 0.9370 ;
      RECT 2.4830 0.6020 2.5330 0.8870 ;
      RECT 1.5500 1.0010 2.6490 1.0510 ;
      RECT 2.5990 0.4960 2.6490 1.0010 ;
      RECT 2.5590 1.0510 2.6090 1.3080 ;
      RECT 2.4070 0.4460 2.6490 0.4960 ;
      RECT 2.4070 1.3080 2.6090 1.3580 ;
      RECT 2.5590 0.3710 2.6090 0.4460 ;
      RECT 2.4070 0.3710 2.4570 0.4460 ;
      RECT 2.4070 1.2160 2.4570 1.3080 ;
      RECT 2.0860 1.1660 2.4570 1.2160 ;
      RECT 3.2070 0.6040 4.2210 0.6540 ;
      RECT 3.2070 0.6540 3.2570 0.9780 ;
      RECT 2.8460 0.9780 3.2570 1.0280 ;
      RECT 2.8460 0.5880 2.8960 0.9780 ;
      RECT 2.8460 0.5380 2.9530 0.5880 ;
      RECT 3.2260 1.4080 3.7650 1.4580 ;
      RECT 1.4190 1.4780 1.9410 1.5280 ;
      RECT 1.4190 1.5280 1.4690 1.5650 ;
      RECT 0.7950 1.5260 1.3170 1.5760 ;
      RECT 1.2670 1.4280 1.3170 1.5260 ;
      RECT 1.2670 1.3780 2.0770 1.4280 ;
      RECT 2.0270 1.4280 2.0770 1.5440 ;
      RECT 0.5830 0.6180 1.0290 0.6680 ;
      RECT 0.5830 0.6680 0.6330 0.9140 ;
      RECT 0.5830 0.4220 0.6330 0.6180 ;
      RECT 1.0390 0.5180 1.1650 0.5680 ;
      RECT 1.0390 0.3940 1.0890 0.5180 ;
      RECT 1.1150 0.5680 1.1650 0.7180 ;
      RECT 1.0390 0.7180 1.1650 0.7680 ;
      RECT 1.0390 0.7680 1.0890 0.9140 ;
      RECT 3.3450 0.7090 3.7650 0.7590 ;
      RECT 3.3450 0.7590 3.3950 1.0990 ;
      RECT 2.8350 1.0990 3.3950 1.1490 ;
      RECT 2.8350 1.1490 2.8850 1.2720 ;
      RECT 2.6590 1.2720 2.8850 1.3220 ;
      RECT 2.6590 1.3220 2.7090 1.4280 ;
      RECT 2.4670 1.4280 2.7090 1.4780 ;
      RECT 1.0990 0.0960 1.4910 0.1460 ;
      RECT 2.2860 1.5280 3.6260 1.5780 ;
      RECT 3.3030 1.2080 3.6890 1.2580 ;
      RECT 1.4790 1.2780 1.8650 1.3280 ;
    LAYER PO ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 1.2770 0.0680 1.3070 0.5420 ;
      RECT 4.3170 0.0680 4.3470 1.6060 ;
      RECT 3.7090 0.0680 3.7390 0.7870 ;
      RECT 2.6450 0.0680 2.6750 0.6220 ;
      RECT 1.8850 0.8530 1.9150 1.6060 ;
      RECT 1.8850 0.0680 1.9150 0.6610 ;
      RECT 2.6450 0.7320 2.6750 1.6060 ;
      RECT 4.4690 0.0680 4.4990 1.6060 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 3.7090 1.0120 3.7390 1.6060 ;
      RECT 1.2770 0.7900 1.3070 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
  END
END DFFNASRQX2_LVT

MACRO DFFNASRX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.56 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.5600 0.0300 ;
        RECT 0.5860 0.0300 0.6360 0.1960 ;
        RECT 0.2790 0.0300 0.3290 0.4190 ;
        RECT 4.0790 0.0300 4.1290 0.2200 ;
        RECT 1.5410 0.0300 1.5910 0.2870 ;
        RECT 3.7750 0.0300 3.8250 0.3300 ;
        RECT 0.5860 0.1960 0.9370 0.2460 ;
        RECT 1.5410 0.2870 2.1530 0.3370 ;
        RECT 3.1510 0.3300 3.8410 0.3800 ;
        RECT 0.8870 0.2460 0.9370 0.4500 ;
        RECT 0.7350 0.2460 0.7850 0.4500 ;
        RECT 2.1030 0.3370 2.1530 0.4610 ;
        RECT 1.9510 0.3370 2.0010 0.4610 ;
    END
  END VSS

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.3530 1.1610 4.4640 1.2210 ;
        RECT 4.2310 1.2210 4.4640 1.2710 ;
        RECT 4.4130 0.2040 4.4630 1.1610 ;
        RECT 4.2310 1.2710 4.2810 1.5460 ;
        RECT 4.2150 0.1540 4.4630 0.2040 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.5600 1.7020 ;
        RECT 0.2790 1.0330 0.3290 1.6420 ;
        RECT 4.0790 0.9470 4.1290 1.6420 ;
        RECT 2.1270 1.3280 2.1770 1.6420 ;
        RECT 3.8150 1.3580 3.8650 1.6420 ;
        RECT 0.4330 1.3580 0.4830 1.6420 ;
        RECT 1.9340 1.2780 2.3360 1.3280 ;
        RECT 2.9860 1.3080 3.8650 1.3580 ;
        RECT 0.4330 1.3380 0.9370 1.3580 ;
        RECT 0.4340 1.3080 0.9370 1.3380 ;
        RECT 0.7350 1.0920 0.7850 1.3080 ;
        RECT 0.8870 1.1050 0.9370 1.3080 ;
    END
  END VDD

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9230 0.1380 3.0050 0.1740 ;
        RECT 1.7230 0.0880 3.0050 0.1380 ;
        RECT 1.7230 0.1380 1.8790 0.2070 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.3590 0.6800 ;
        RECT 0.2490 0.6800 0.4210 0.7300 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.5310 0.8570 3.7030 1.0340 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.4240 0.7250 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.2010 1.0090 4.3110 1.1190 ;
        RECT 4.2610 0.8540 4.3110 1.0090 ;
        RECT 3.9270 0.8040 4.3110 0.8540 ;
        RECT 3.9270 0.8540 3.9770 1.5460 ;
        RECT 4.2610 0.3590 4.3110 0.8040 ;
        RECT 3.9270 0.3090 4.3110 0.3590 ;
        RECT 3.9270 0.1480 3.9770 0.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 4.6750 1.7730 ;
    LAYER M1 ;
      RECT 1.8590 0.8820 2.5330 0.9320 ;
      RECT 2.4830 0.5970 2.5330 0.8820 ;
      RECT 1.1910 0.2990 1.2810 0.3810 ;
      RECT 1.2150 0.3810 1.2650 0.9880 ;
      RECT 0.4310 0.9880 1.2650 1.0380 ;
      RECT 1.1910 1.0380 1.2410 1.3140 ;
      RECT 0.4310 1.0380 0.4810 1.2160 ;
      RECT 0.4310 0.8290 0.4810 0.9880 ;
      RECT 0.4310 0.5790 0.5210 0.6290 ;
      RECT 0.4310 0.4550 0.4810 0.5790 ;
      RECT 0.4310 0.7800 0.5210 0.8290 ;
      RECT 0.4710 0.6290 0.5210 0.7800 ;
      RECT 3.2430 0.0880 3.2930 0.2300 ;
      RECT 2.2950 0.2300 3.2930 0.2800 ;
      RECT 2.6190 0.2800 2.7010 0.3000 ;
      RECT 2.6190 0.1980 2.7010 0.2300 ;
      RECT 2.2950 0.2800 2.3450 0.5840 ;
      RECT 1.8590 0.5840 2.3450 0.6340 ;
      RECT 1.3430 0.6840 2.2450 0.7340 ;
      RECT 1.3430 0.7340 1.3930 1.1580 ;
      RECT 1.3430 0.4840 1.3930 0.6840 ;
      RECT 1.3430 1.2080 1.3930 1.3140 ;
      RECT 1.3430 0.3550 1.3930 0.4340 ;
      RECT 1.3430 1.1580 1.7130 1.2080 ;
      RECT 1.3430 0.4340 1.5610 0.4840 ;
      RECT 4.1550 0.4880 4.2050 0.7040 ;
      RECT 2.7110 0.4380 4.2050 0.4880 ;
      RECT 3.8150 0.7040 4.2050 0.7540 ;
      RECT 3.8150 0.7540 3.8650 1.1080 ;
      RECT 3.4550 1.1080 3.8650 1.1580 ;
      RECT 2.7110 0.4880 2.7610 1.1650 ;
      RECT 3.0140 0.4880 3.0640 0.7660 ;
      RECT 3.0140 0.7660 3.1570 0.8160 ;
      RECT 1.5500 1.0010 2.6490 1.0510 ;
      RECT 2.5990 0.4960 2.6490 1.0010 ;
      RECT 2.5590 1.0510 2.6090 1.3080 ;
      RECT 2.4070 0.4460 2.6490 0.4960 ;
      RECT 2.4070 1.3080 2.6090 1.3580 ;
      RECT 2.5590 0.3710 2.6090 0.4460 ;
      RECT 2.4070 0.3710 2.4570 0.4460 ;
      RECT 2.4070 1.2160 2.4570 1.3080 ;
      RECT 2.0860 1.1660 2.4570 1.2160 ;
      RECT 3.2070 0.6040 4.0690 0.6540 ;
      RECT 3.2070 0.6540 3.2570 0.9780 ;
      RECT 2.8460 0.9780 3.2570 1.0280 ;
      RECT 2.8460 0.5880 2.8960 0.9780 ;
      RECT 2.8460 0.5380 2.9530 0.5880 ;
      RECT 3.2260 1.4080 3.7650 1.4580 ;
      RECT 1.4190 1.4780 1.9410 1.5280 ;
      RECT 1.4190 1.5280 1.4690 1.5650 ;
      RECT 0.7950 1.5260 1.3170 1.5760 ;
      RECT 1.2670 1.4280 1.3170 1.5260 ;
      RECT 1.2670 1.3780 2.0770 1.4280 ;
      RECT 2.0270 1.4280 2.0770 1.5440 ;
      RECT 0.5830 0.6180 1.0290 0.6680 ;
      RECT 0.5830 0.6680 0.6330 0.9140 ;
      RECT 0.5830 0.4220 0.6330 0.6180 ;
      RECT 1.0390 0.5180 1.1650 0.5680 ;
      RECT 1.0390 0.3940 1.0890 0.5180 ;
      RECT 1.1150 0.5680 1.1650 0.7180 ;
      RECT 1.0390 0.7180 1.1650 0.7680 ;
      RECT 1.0390 0.7680 1.0890 0.9140 ;
      RECT 3.3450 0.7090 3.7650 0.7590 ;
      RECT 3.3450 0.7590 3.3950 1.0990 ;
      RECT 2.8350 1.0990 3.3950 1.1490 ;
      RECT 2.8350 1.1490 2.8850 1.2720 ;
      RECT 2.6590 1.2720 2.8850 1.3220 ;
      RECT 2.6590 1.3220 2.7090 1.4280 ;
      RECT 2.4670 1.4280 2.7090 1.4780 ;
      RECT 1.0990 0.0960 1.4910 0.1460 ;
      RECT 2.2860 1.5280 3.6260 1.5780 ;
      RECT 3.3030 1.2080 3.6890 1.2580 ;
      RECT 1.4790 1.2780 1.8650 1.3280 ;
    LAYER PO ;
      RECT 4.3170 0.0680 4.3470 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 1.2770 0.0680 1.3070 0.5420 ;
      RECT 4.4690 0.0680 4.4990 1.6060 ;
      RECT 1.2770 0.7900 1.3070 1.6060 ;
      RECT 3.7090 0.0680 3.7390 0.7870 ;
      RECT 1.8850 0.0680 1.9150 0.6620 ;
      RECT 3.7090 1.0120 3.7390 1.6060 ;
      RECT 2.6450 0.7320 2.6750 1.6060 ;
      RECT 2.6450 0.0680 2.6750 0.6220 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 1.8850 0.8540 1.9150 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
  END
END DFFNASRX1_LVT

MACRO DFFNASRX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.864 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6570 0.2170 4.7670 0.2700 ;
        RECT 4.3830 0.2700 4.7670 0.3200 ;
        RECT 4.6570 0.3200 4.7670 0.3590 ;
        RECT 4.3830 0.1480 4.4330 0.2700 ;
        RECT 4.6990 0.3590 4.7490 0.9180 ;
        RECT 4.3830 0.9180 4.7490 0.9680 ;
        RECT 4.3830 0.9680 4.4330 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.8640 0.0300 ;
        RECT 0.5860 0.0300 0.6360 0.1960 ;
        RECT 3.9270 0.0300 3.9770 0.4080 ;
        RECT 0.2790 0.0300 0.3290 0.4190 ;
        RECT 4.5350 0.0300 4.5850 0.2200 ;
        RECT 4.2320 0.0300 4.2820 0.3120 ;
        RECT 1.5410 0.0300 1.5910 0.2870 ;
        RECT 3.7750 0.0300 3.8250 0.3300 ;
        RECT 0.5860 0.1960 0.9370 0.2460 ;
        RECT 1.5410 0.2870 2.1530 0.3370 ;
        RECT 3.1510 0.3300 3.8410 0.3800 ;
        RECT 0.8870 0.2460 0.9370 0.4500 ;
        RECT 0.7350 0.2460 0.7850 0.4500 ;
        RECT 2.1030 0.3370 2.1530 0.4610 ;
        RECT 1.9510 0.3370 2.0010 0.4610 ;
    END
  END VSS

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0790 0.1480 4.1290 0.3940 ;
        RECT 4.0790 0.3940 4.5870 0.4010 ;
        RECT 4.0790 0.4010 4.6250 0.4440 ;
        RECT 4.5050 0.4440 4.6250 0.5110 ;
        RECT 4.5750 0.5110 4.6250 0.8040 ;
        RECT 4.0790 0.8040 4.6250 0.8540 ;
        RECT 4.0790 0.8540 4.1290 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.8640 1.7020 ;
        RECT 0.2790 1.0330 0.3290 1.6420 ;
        RECT 4.2310 0.9600 4.2810 1.6420 ;
        RECT 3.9270 0.9120 3.9770 1.6420 ;
        RECT 4.5350 1.0520 4.5850 1.6420 ;
        RECT 2.1270 1.3280 2.1770 1.6420 ;
        RECT 3.8150 1.3580 3.8650 1.6420 ;
        RECT 0.4330 1.3580 0.4830 1.6420 ;
        RECT 1.9340 1.2780 2.3360 1.3280 ;
        RECT 2.9860 1.3080 3.8650 1.3580 ;
        RECT 0.4330 1.3380 0.9370 1.3580 ;
        RECT 0.4340 1.3080 0.9370 1.3380 ;
        RECT 0.7350 1.0920 0.7850 1.3080 ;
        RECT 0.8870 1.1050 0.9370 1.3080 ;
    END
  END VDD

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7230 0.0900 3.0050 0.1400 ;
        RECT 2.9230 0.1400 3.0050 0.1760 ;
        RECT 1.7230 0.1400 1.8790 0.2190 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END RSTB

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.3590 0.6800 ;
        RECT 0.2490 0.6800 0.4210 0.7300 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.5310 0.8570 3.7030 1.0340 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.4240 0.7250 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 4.9790 1.7730 ;
    LAYER M1 ;
      RECT 4.2880 0.6040 4.5250 0.6540 ;
      RECT 3.8150 0.7540 3.8650 1.1080 ;
      RECT 3.4550 1.1080 3.8650 1.1580 ;
      RECT 4.2880 0.5460 4.3380 0.6040 ;
      RECT 4.2880 0.6540 4.3380 0.7040 ;
      RECT 3.0140 0.4960 4.3380 0.5460 ;
      RECT 3.8150 0.7040 4.3380 0.7540 ;
      RECT 3.0140 0.4880 3.0640 0.4960 ;
      RECT 3.0140 0.5460 3.0640 0.7660 ;
      RECT 2.7110 0.4380 3.0640 0.4880 ;
      RECT 3.0140 0.7660 3.1570 0.8160 ;
      RECT 2.7110 0.4880 2.7610 1.1650 ;
      RECT 1.8590 0.8820 2.5330 0.9320 ;
      RECT 2.4830 0.5970 2.5330 0.8820 ;
      RECT 1.1910 0.2990 1.2810 0.3810 ;
      RECT 1.2150 0.3810 1.2650 0.9880 ;
      RECT 0.4310 0.9880 1.2650 1.0380 ;
      RECT 1.1910 1.0380 1.2410 1.3140 ;
      RECT 0.4310 1.0380 0.4810 1.2160 ;
      RECT 0.4310 0.8290 0.4810 0.9880 ;
      RECT 0.4310 0.5790 0.5210 0.6290 ;
      RECT 0.4310 0.4550 0.4810 0.5790 ;
      RECT 0.4310 0.7800 0.5210 0.8290 ;
      RECT 0.4710 0.6290 0.5210 0.7800 ;
      RECT 3.2430 0.1020 3.2930 0.2300 ;
      RECT 2.2950 0.2300 3.2930 0.2800 ;
      RECT 2.6190 0.1980 2.7010 0.2300 ;
      RECT 2.2950 0.2800 2.3450 0.5840 ;
      RECT 1.8590 0.5840 2.3450 0.6340 ;
      RECT 1.3430 0.6840 2.2450 0.7340 ;
      RECT 1.3430 0.7340 1.3930 1.1580 ;
      RECT 1.3430 0.4840 1.3930 0.6840 ;
      RECT 1.3430 1.2080 1.3930 1.3140 ;
      RECT 1.3430 0.3550 1.3930 0.4340 ;
      RECT 1.3430 1.1580 1.7130 1.2080 ;
      RECT 1.3430 0.4340 1.5610 0.4840 ;
      RECT 1.5500 1.0010 2.6490 1.0510 ;
      RECT 2.5990 0.4960 2.6490 1.0010 ;
      RECT 2.5590 1.0510 2.6090 1.3080 ;
      RECT 2.4070 0.4460 2.6490 0.4960 ;
      RECT 2.4070 1.3080 2.6090 1.3580 ;
      RECT 2.5590 0.3710 2.6090 0.4460 ;
      RECT 2.4070 0.3710 2.4570 0.4460 ;
      RECT 2.4070 1.2160 2.4570 1.3080 ;
      RECT 2.0860 1.1660 2.4570 1.2160 ;
      RECT 3.2070 0.6040 4.2210 0.6540 ;
      RECT 3.2070 0.6540 3.2570 0.9780 ;
      RECT 2.8460 0.9780 3.2570 1.0280 ;
      RECT 2.8460 0.5880 2.8960 0.9780 ;
      RECT 2.8460 0.5380 2.9530 0.5880 ;
      RECT 3.2260 1.4080 3.7650 1.4580 ;
      RECT 1.4190 1.4780 1.9410 1.5280 ;
      RECT 1.4190 1.5280 1.4690 1.5650 ;
      RECT 0.7950 1.5260 1.3170 1.5760 ;
      RECT 1.2670 1.4280 1.3170 1.5260 ;
      RECT 1.2670 1.3780 2.0770 1.4280 ;
      RECT 2.0270 1.4280 2.0770 1.5440 ;
      RECT 0.5830 0.6180 1.0290 0.6680 ;
      RECT 0.5830 0.6680 0.6330 0.9140 ;
      RECT 0.5830 0.4220 0.6330 0.6180 ;
      RECT 1.0390 0.5180 1.1650 0.5680 ;
      RECT 1.0390 0.3940 1.0890 0.5180 ;
      RECT 1.1150 0.5680 1.1650 0.7180 ;
      RECT 1.0390 0.7180 1.1650 0.7680 ;
      RECT 1.0390 0.7680 1.0890 0.9140 ;
      RECT 3.3450 0.7090 3.7650 0.7590 ;
      RECT 3.3450 0.7590 3.3950 1.0990 ;
      RECT 2.8350 1.0990 3.3950 1.1490 ;
      RECT 2.8350 1.1490 2.8850 1.2720 ;
      RECT 2.6590 1.2720 2.8850 1.3220 ;
      RECT 2.6590 1.3220 2.7090 1.4280 ;
      RECT 2.4670 1.4280 2.7090 1.4780 ;
      RECT 1.0990 0.0960 1.4910 0.1460 ;
      RECT 2.2860 1.5280 3.6260 1.5780 ;
      RECT 3.3030 1.2080 3.6890 1.2580 ;
      RECT 1.4790 1.2780 1.8650 1.3280 ;
    LAYER PO ;
      RECT 3.7090 1.0120 3.7390 1.6060 ;
      RECT 2.6450 0.7320 2.6750 1.6060 ;
      RECT 2.6450 0.0680 2.6750 0.6220 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 1.8850 0.8540 1.9150 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 4.6210 0.0680 4.6510 1.6060 ;
      RECT 1.2770 0.0680 1.3070 0.5420 ;
      RECT 1.2770 0.7900 1.3070 1.6060 ;
      RECT 4.7730 0.0680 4.8030 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 4.4690 0.0680 4.4990 1.6060 ;
      RECT 3.7090 0.0680 3.7390 0.7870 ;
      RECT 1.8850 0.0680 1.9150 0.6620 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 4.3170 0.0680 4.3470 1.6060 ;
  END
END DFFNASRX2_LVT

MACRO DFFNASX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.256 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.2560 0.0300 ;
        RECT 0.5860 0.0300 0.6360 0.1960 ;
        RECT 0.2790 0.0300 0.3290 0.4190 ;
        RECT 1.9510 0.0300 2.0010 0.4610 ;
        RECT 3.7750 0.0300 3.8250 0.2200 ;
        RECT 3.4710 0.0300 3.5210 0.3300 ;
        RECT 1.7990 0.0300 1.8490 0.3710 ;
        RECT 0.5860 0.1960 0.9370 0.2460 ;
        RECT 2.8450 0.3300 3.5370 0.3800 ;
        RECT 0.8870 0.2460 0.9370 0.4500 ;
        RECT 0.7350 0.2460 0.7850 0.4500 ;
    END
  END VSS

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0490 1.1610 4.1600 1.2210 ;
        RECT 3.9270 1.2210 4.1600 1.2710 ;
        RECT 4.1090 0.2040 4.1590 1.1610 ;
        RECT 3.9270 1.2710 3.9770 1.5460 ;
        RECT 3.9110 0.1540 4.1590 0.2040 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.2560 1.7020 ;
        RECT 0.2790 1.0330 0.3290 1.6420 ;
        RECT 3.7750 0.9470 3.8250 1.6420 ;
        RECT 1.9750 1.3210 2.0250 1.6420 ;
        RECT 3.5110 1.3580 3.5610 1.6420 ;
        RECT 0.4330 1.3600 0.4830 1.6420 ;
        RECT 1.7740 1.2710 2.1840 1.3210 ;
        RECT 2.8340 1.3080 3.5610 1.3580 ;
        RECT 0.4330 1.3400 0.9370 1.3600 ;
        RECT 0.4340 1.3100 0.9370 1.3400 ;
        RECT 0.7350 1.0940 0.7850 1.3100 ;
        RECT 0.8870 1.1070 0.9370 1.3100 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.3590 0.6800 ;
        RECT 0.2490 0.6800 0.4210 0.7300 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2270 0.8570 3.3990 1.0340 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.4240 0.7250 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8970 1.0090 4.0070 1.1190 ;
        RECT 3.9570 0.8540 4.0070 1.0090 ;
        RECT 3.6230 0.8040 4.0070 0.8540 ;
        RECT 3.6230 0.8540 3.6730 1.5460 ;
        RECT 3.9570 0.3590 4.0070 0.8040 ;
        RECT 3.6230 0.3090 4.0070 0.3590 ;
        RECT 3.6230 0.1480 3.6730 0.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 4.3710 1.7730 ;
    LAYER M1 ;
      RECT 1.1910 0.2990 1.2810 0.3810 ;
      RECT 1.2150 0.3810 1.2650 0.9880 ;
      RECT 0.4310 0.9880 1.2650 1.0380 ;
      RECT 1.1910 1.0380 1.2410 1.3140 ;
      RECT 0.4310 1.0380 0.4810 1.2160 ;
      RECT 0.4310 0.8290 0.4810 0.9880 ;
      RECT 0.4310 0.5790 0.5210 0.6290 ;
      RECT 0.4310 0.4550 0.4810 0.5790 ;
      RECT 0.4310 0.7800 0.5210 0.8290 ;
      RECT 0.4710 0.6290 0.5210 0.7800 ;
      RECT 2.9390 0.0880 2.9890 0.2300 ;
      RECT 2.1430 0.2300 2.9890 0.2800 ;
      RECT 2.4670 0.1780 2.5490 0.2300 ;
      RECT 2.1430 0.2800 2.1930 0.5840 ;
      RECT 1.7060 0.5840 2.1930 0.6340 ;
      RECT 2.1430 0.6340 2.1930 0.6360 ;
      RECT 3.8510 0.4810 3.9010 0.7040 ;
      RECT 2.5590 0.4310 3.9010 0.4810 ;
      RECT 3.5110 0.7040 3.9010 0.7540 ;
      RECT 3.5110 0.7540 3.5610 1.1080 ;
      RECT 3.1510 1.1080 3.5610 1.1580 ;
      RECT 2.5590 0.4810 2.6090 1.1650 ;
      RECT 2.8270 0.4810 2.8770 0.6960 ;
      RECT 2.7710 0.6960 2.8770 0.7460 ;
      RECT 1.6980 0.8780 2.3810 0.9280 ;
      RECT 2.3310 0.5970 2.3810 0.8780 ;
      RECT 1.3430 0.7440 2.0930 0.7940 ;
      RECT 1.3430 0.7940 1.3930 1.1560 ;
      RECT 1.3430 0.4820 1.3930 0.7440 ;
      RECT 1.3430 1.1560 1.5610 1.2060 ;
      RECT 1.3430 0.4320 1.5610 0.4820 ;
      RECT 1.3430 1.2060 1.3930 1.3140 ;
      RECT 1.3430 0.3550 1.3930 0.4320 ;
      RECT 1.4190 1.4760 1.7890 1.5260 ;
      RECT 1.4190 1.5260 1.4690 1.5630 ;
      RECT 2.9530 0.6040 3.7650 0.6050 ;
      RECT 2.9320 0.6050 3.7650 0.6540 ;
      RECT 2.9320 0.6540 2.9820 0.9750 ;
      RECT 2.6710 0.9750 2.9820 1.0240 ;
      RECT 2.6880 1.0240 2.9820 1.0250 ;
      RECT 2.6710 0.5850 2.7210 0.9750 ;
      RECT 2.6710 0.5350 2.7770 0.5850 ;
      RECT 3.0510 0.7090 3.4610 0.7590 ;
      RECT 3.0510 0.7590 3.1010 1.0990 ;
      RECT 2.6830 1.0990 3.1010 1.1490 ;
      RECT 2.6830 1.1490 2.7330 1.2720 ;
      RECT 2.6830 1.0960 2.7330 1.0990 ;
      RECT 2.5070 1.2720 2.7330 1.3220 ;
      RECT 2.5070 1.3220 2.5570 1.4280 ;
      RECT 2.3150 1.4280 2.5570 1.4780 ;
      RECT 1.5500 1.0010 2.4970 1.0510 ;
      RECT 2.4470 0.4960 2.4970 1.0010 ;
      RECT 2.4070 1.0510 2.4570 1.3080 ;
      RECT 2.2550 0.4460 2.4970 0.4960 ;
      RECT 2.2550 1.3080 2.4570 1.3580 ;
      RECT 2.4070 0.3710 2.4570 0.4460 ;
      RECT 2.2550 0.3710 2.3050 0.4460 ;
      RECT 2.2550 1.2160 2.3050 1.3080 ;
      RECT 1.9340 1.1660 2.3050 1.2160 ;
      RECT 0.7950 1.5260 1.3170 1.5760 ;
      RECT 1.2670 1.4260 1.3170 1.5260 ;
      RECT 1.2670 1.3760 1.9250 1.4260 ;
      RECT 1.8750 1.4260 1.9250 1.5840 ;
      RECT 2.9220 1.5190 3.4610 1.5690 ;
      RECT 0.5830 0.6180 1.0290 0.6680 ;
      RECT 0.5830 0.6680 0.6330 0.9140 ;
      RECT 0.5830 0.4220 0.6330 0.6180 ;
      RECT 1.0390 0.5180 1.1650 0.5680 ;
      RECT 1.0390 0.3940 1.0890 0.5180 ;
      RECT 1.1150 0.5680 1.1650 0.7180 ;
      RECT 1.0390 0.7180 1.1650 0.7680 ;
      RECT 1.0390 0.7680 1.0890 0.9140 ;
      RECT 2.1340 1.5280 2.6820 1.5780 ;
      RECT 2.6320 1.4610 2.6820 1.5280 ;
      RECT 2.6320 1.4110 3.3090 1.4610 ;
      RECT 1.0990 0.0960 1.4910 0.1460 ;
      RECT 2.9990 1.2080 3.3850 1.2580 ;
    LAYER PO ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 3.7090 0.0680 3.7390 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 2.4930 0.7270 2.5230 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 1.2770 0.0680 1.3070 0.5420 ;
      RECT 1.8850 0.0660 1.9150 1.6040 ;
      RECT 3.4050 0.0680 3.4350 0.7870 ;
      RECT 2.7970 0.0650 2.8270 1.6030 ;
      RECT 1.5810 0.0660 1.6110 1.6040 ;
      RECT 1.4290 0.0660 1.4590 1.6040 ;
      RECT 1.7330 0.0660 1.7630 0.6620 ;
      RECT 1.2770 0.7900 1.3070 1.6060 ;
      RECT 3.4050 1.0120 3.4350 1.6060 ;
      RECT 1.7330 0.8300 1.7630 1.6040 ;
      RECT 2.4930 0.0680 2.5230 0.6220 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
  END
END DFFNASX1_LVT

MACRO DFFNASX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.56 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.3530 0.0970 4.4630 0.2070 ;
        RECT 4.3950 0.2070 4.4450 0.2700 ;
        RECT 4.0790 0.2700 4.4450 0.3200 ;
        RECT 4.0790 0.1480 4.1290 0.2700 ;
        RECT 4.3950 0.3200 4.4450 0.9180 ;
        RECT 4.0790 0.9180 4.4450 0.9680 ;
        RECT 4.0790 0.9680 4.1290 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.7750 0.1480 3.8250 0.3940 ;
        RECT 3.7750 0.3940 4.3210 0.4440 ;
        RECT 4.2010 0.4440 4.3210 0.5110 ;
        RECT 4.2710 0.5110 4.3210 0.8040 ;
        RECT 3.7750 0.8040 4.3210 0.8540 ;
        RECT 3.7750 0.8540 3.8250 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.5600 0.0300 ;
        RECT 0.5860 0.0300 0.6360 0.1960 ;
        RECT 4.2310 0.0300 4.2810 0.2200 ;
        RECT 3.9280 0.0300 3.9780 0.3120 ;
        RECT 3.6230 0.0300 3.6730 0.4080 ;
        RECT 0.2790 0.0300 0.3290 0.4190 ;
        RECT 1.9510 0.0300 2.0010 0.4610 ;
        RECT 1.7990 0.0300 1.8490 0.3710 ;
        RECT 3.4710 0.0300 3.5210 0.3300 ;
        RECT 0.5860 0.1960 0.9370 0.2460 ;
        RECT 2.8450 0.3300 3.5370 0.3800 ;
        RECT 0.8870 0.2460 0.9370 0.4500 ;
        RECT 0.7350 0.2460 0.7850 0.4500 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.5600 1.7020 ;
        RECT 0.2790 1.0330 0.3290 1.6420 ;
        RECT 3.6230 0.9120 3.6730 1.6420 ;
        RECT 3.9270 0.9600 3.9770 1.6420 ;
        RECT 4.2310 1.0520 4.2810 1.6420 ;
        RECT 1.9750 1.3210 2.0250 1.6420 ;
        RECT 3.5110 1.3580 3.5610 1.6420 ;
        RECT 0.4330 1.3600 0.4830 1.6420 ;
        RECT 1.7740 1.2710 2.1840 1.3210 ;
        RECT 2.8340 1.3080 3.5610 1.3580 ;
        RECT 0.4330 1.3400 0.9370 1.3600 ;
        RECT 0.4340 1.3100 0.9370 1.3400 ;
        RECT 0.7350 1.0940 0.7850 1.3100 ;
        RECT 0.8870 1.1070 0.9370 1.3100 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.3590 0.6800 ;
        RECT 0.2490 0.6800 0.4210 0.7300 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2270 0.8570 3.3990 1.0340 ;
    END
    ANTENNAGATEAREA 0.042 ;
  END SETB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.4240 0.7250 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 4.6750 1.7730 ;
    LAYER M1 ;
      RECT 1.1910 0.2990 1.2810 0.3810 ;
      RECT 1.2150 0.3810 1.2650 0.9880 ;
      RECT 0.4310 0.9880 1.2650 1.0380 ;
      RECT 1.1910 1.0380 1.2410 1.3140 ;
      RECT 0.4310 1.0380 0.4810 1.2160 ;
      RECT 0.4310 0.8290 0.4810 0.9880 ;
      RECT 0.4310 0.5790 0.5210 0.6290 ;
      RECT 0.4310 0.4550 0.4810 0.5790 ;
      RECT 0.4310 0.7800 0.5210 0.8290 ;
      RECT 0.4710 0.6290 0.5210 0.7800 ;
      RECT 2.9390 0.0880 2.9890 0.2300 ;
      RECT 2.1430 0.2300 2.9890 0.2800 ;
      RECT 2.4670 0.1780 2.5490 0.2300 ;
      RECT 2.1430 0.2800 2.1930 0.5840 ;
      RECT 1.7060 0.5840 2.1930 0.6340 ;
      RECT 2.1430 0.6340 2.1930 0.6360 ;
      RECT 3.9840 0.6040 4.2210 0.6540 ;
      RECT 3.5110 0.7540 3.5610 1.1080 ;
      RECT 3.1510 1.1080 3.5610 1.1580 ;
      RECT 3.9840 0.6540 4.0340 0.7040 ;
      RECT 3.9840 0.5490 4.0340 0.6040 ;
      RECT 2.8270 0.4990 4.0340 0.5490 ;
      RECT 3.5110 0.7040 4.0340 0.7540 ;
      RECT 2.8270 0.5490 2.8770 0.6960 ;
      RECT 2.8270 0.4810 2.8770 0.4990 ;
      RECT 2.7710 0.6960 2.8770 0.7460 ;
      RECT 2.5590 0.4310 2.8770 0.4810 ;
      RECT 2.5590 0.4810 2.6090 1.1650 ;
      RECT 1.6980 0.8780 2.3810 0.9280 ;
      RECT 2.3310 0.5970 2.3810 0.8780 ;
      RECT 1.3430 0.7440 2.0930 0.7940 ;
      RECT 1.3430 0.7940 1.3930 1.1560 ;
      RECT 1.3430 0.4820 1.3930 0.7440 ;
      RECT 1.3430 1.1560 1.5610 1.2060 ;
      RECT 1.3430 0.4320 1.5610 0.4820 ;
      RECT 1.3430 1.2060 1.3930 1.3140 ;
      RECT 1.3430 0.3550 1.3930 0.4320 ;
      RECT 1.5500 1.0010 2.4970 1.0510 ;
      RECT 2.4070 1.0510 2.4570 1.3080 ;
      RECT 2.4470 0.4960 2.4970 1.0010 ;
      RECT 2.2550 1.3080 2.4570 1.3580 ;
      RECT 2.2550 0.4460 2.4970 0.4960 ;
      RECT 2.2550 1.2160 2.3050 1.3080 ;
      RECT 2.4070 0.3710 2.4570 0.4460 ;
      RECT 2.2550 0.3710 2.3050 0.4460 ;
      RECT 1.9340 1.1660 2.3050 1.2160 ;
      RECT 2.9530 0.6040 3.9170 0.6050 ;
      RECT 2.9320 0.6050 3.9170 0.6540 ;
      RECT 2.9320 0.6540 2.9820 0.9750 ;
      RECT 2.6710 0.9750 2.9820 1.0240 ;
      RECT 2.6710 0.5850 2.7210 0.9750 ;
      RECT 2.6880 1.0240 2.9820 1.0250 ;
      RECT 2.6710 0.5350 2.7770 0.5850 ;
      RECT 1.4190 1.4760 1.7890 1.5260 ;
      RECT 1.4190 1.5260 1.4690 1.5630 ;
      RECT 3.0510 0.7090 3.4610 0.7590 ;
      RECT 3.0510 0.7590 3.1010 1.0990 ;
      RECT 2.6830 1.0990 3.1010 1.1490 ;
      RECT 2.6830 1.1490 2.7330 1.2720 ;
      RECT 2.6830 1.0960 2.7330 1.0990 ;
      RECT 2.5070 1.2720 2.7330 1.3220 ;
      RECT 2.5070 1.3220 2.5570 1.4280 ;
      RECT 2.3150 1.4280 2.5570 1.4780 ;
      RECT 0.7950 1.5260 1.3170 1.5760 ;
      RECT 1.2670 1.4260 1.3170 1.5260 ;
      RECT 1.2670 1.3760 1.9250 1.4260 ;
      RECT 1.8750 1.4260 1.9250 1.5840 ;
      RECT 2.9220 1.5190 3.4610 1.5690 ;
      RECT 0.5830 0.6180 1.0290 0.6680 ;
      RECT 0.5830 0.6680 0.6330 0.9140 ;
      RECT 0.5830 0.4220 0.6330 0.6180 ;
      RECT 1.0390 0.5180 1.1650 0.5680 ;
      RECT 1.0390 0.3940 1.0890 0.5180 ;
      RECT 1.1150 0.5680 1.1650 0.7180 ;
      RECT 1.0390 0.7180 1.1650 0.7680 ;
      RECT 1.0390 0.7680 1.0890 0.9140 ;
      RECT 2.1340 1.5280 2.6820 1.5780 ;
      RECT 2.6320 1.4610 2.6820 1.5280 ;
      RECT 2.6320 1.4110 3.3090 1.4610 ;
      RECT 1.0990 0.0960 1.4910 0.1460 ;
      RECT 2.9990 1.2080 3.3850 1.2580 ;
    LAYER PO ;
      RECT 1.7330 0.8300 1.7630 1.6040 ;
      RECT 2.4930 0.0680 2.5230 0.6220 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 2.4930 0.7270 2.5230 1.6060 ;
      RECT 4.3170 0.0680 4.3470 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 4.4690 0.0680 4.4990 1.6060 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 3.7090 0.0680 3.7390 1.6060 ;
      RECT 1.2770 0.0680 1.3070 0.5420 ;
      RECT 1.8850 0.0660 1.9150 1.6040 ;
      RECT 3.4050 0.0680 3.4350 0.7870 ;
      RECT 2.7970 0.0650 2.8270 1.6030 ;
      RECT 1.5810 0.0660 1.6110 1.6040 ;
      RECT 1.4290 0.0660 1.4590 1.6040 ;
      RECT 1.7330 0.0660 1.7630 0.6620 ;
      RECT 1.2770 0.7900 1.3070 1.6060 ;
      RECT 3.4050 1.0120 3.4350 1.6060 ;
  END
END DFFNASX2_LVT

MACRO DFFNX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.952 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.9520 0.0300 ;
        RECT 0.5860 0.0300 0.6360 0.1960 ;
        RECT 1.7990 0.0300 1.8490 0.1990 ;
        RECT 0.2790 0.0300 0.3290 0.4190 ;
        RECT 3.4710 0.0300 3.5210 0.2200 ;
        RECT 3.1670 0.0300 3.2170 0.3300 ;
        RECT 0.5860 0.1960 0.9370 0.2460 ;
        RECT 1.7990 0.1990 2.0240 0.2490 ;
        RECT 2.6950 0.3300 3.2330 0.3800 ;
        RECT 0.8870 0.2460 0.9370 0.4500 ;
        RECT 0.7350 0.2460 0.7850 0.4500 ;
        RECT 1.7990 0.2490 1.8490 0.3730 ;
    END
  END VSS

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.7460 1.1610 3.8560 1.2210 ;
        RECT 3.6230 1.2210 3.8560 1.2710 ;
        RECT 3.8050 0.2040 3.8550 1.1610 ;
        RECT 3.6230 1.2710 3.6730 1.5460 ;
        RECT 3.6070 0.1540 3.8550 0.2040 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.9520 1.7020 ;
        RECT 0.2790 1.0330 0.3290 1.6420 ;
        RECT 3.4710 0.9470 3.5210 1.6420 ;
        RECT 2.6390 1.3580 2.6890 1.6420 ;
        RECT 1.9750 1.3280 2.0250 1.6420 ;
        RECT 3.2070 1.3580 3.2570 1.6420 ;
        RECT 0.4330 1.3540 0.4830 1.6420 ;
        RECT 2.6390 1.3080 2.7770 1.3580 ;
        RECT 1.7820 1.2780 2.0250 1.3280 ;
        RECT 3.1490 1.3080 3.2570 1.3580 ;
        RECT 0.4330 1.3340 0.9370 1.3540 ;
        RECT 0.4340 1.3040 0.9370 1.3340 ;
        RECT 0.7350 1.0880 0.7850 1.3040 ;
        RECT 0.8870 1.1010 0.9370 1.3040 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.3590 0.6800 ;
        RECT 0.2490 0.6800 0.4210 0.7300 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.4240 0.7250 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.5930 1.0090 3.7030 1.1190 ;
        RECT 3.6530 0.8540 3.7030 1.0090 ;
        RECT 3.3190 0.8040 3.7030 0.8540 ;
        RECT 3.3190 0.8540 3.3690 1.5460 ;
        RECT 3.6530 0.3590 3.7030 0.8040 ;
        RECT 3.3190 0.3090 3.7030 0.3590 ;
        RECT 3.3190 0.1480 3.3690 0.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 4.0670 1.7730 ;
    LAYER M1 ;
      RECT 1.1910 0.2990 1.2810 0.3810 ;
      RECT 1.2150 0.3810 1.2650 0.9880 ;
      RECT 1.1910 1.0380 1.2410 1.3140 ;
      RECT 0.4310 0.9880 1.2650 1.0380 ;
      RECT 0.4310 1.0380 0.4810 1.2160 ;
      RECT 0.4310 0.8290 0.4810 0.9880 ;
      RECT 0.4310 0.5790 0.5210 0.6290 ;
      RECT 0.4310 0.4550 0.4810 0.5790 ;
      RECT 0.4310 0.7800 0.5210 0.8290 ;
      RECT 0.4710 0.6290 0.5210 0.7800 ;
      RECT 2.7870 0.0880 2.8370 0.2300 ;
      RECT 2.1150 0.2300 2.8370 0.2800 ;
      RECT 2.3150 0.1780 2.3970 0.2300 ;
      RECT 2.1150 0.2800 2.1650 0.3140 ;
      RECT 1.9640 0.3140 2.1650 0.3640 ;
      RECT 1.9640 0.3640 2.0140 0.5400 ;
      RECT 1.7070 0.5400 2.0140 0.5900 ;
      RECT 1.3430 0.6400 2.0930 0.6900 ;
      RECT 1.3430 0.6900 1.3930 1.1580 ;
      RECT 1.3430 0.4840 1.3930 0.6400 ;
      RECT 1.3430 1.1580 1.5610 1.2080 ;
      RECT 1.3430 0.4340 1.5610 0.4840 ;
      RECT 1.3430 1.2080 1.3930 1.3140 ;
      RECT 1.3430 0.3550 1.3930 0.4340 ;
      RECT 3.5470 0.4880 3.5970 0.7040 ;
      RECT 2.4070 0.4380 3.5970 0.4880 ;
      RECT 3.2070 0.7040 3.5970 0.7540 ;
      RECT 3.2070 0.7540 3.2570 1.2080 ;
      RECT 2.8470 1.2080 3.2570 1.2580 ;
      RECT 2.4070 0.4880 2.4570 1.1650 ;
      RECT 2.7100 0.4880 2.7600 0.6990 ;
      RECT 2.6190 0.6990 2.7600 0.7490 ;
      RECT 1.7070 0.7580 2.2290 0.8080 ;
      RECT 2.1790 0.5870 2.2290 0.7580 ;
      RECT 1.5500 1.0010 2.3450 1.0510 ;
      RECT 2.2950 0.4700 2.3450 1.0010 ;
      RECT 2.2550 1.0510 2.3050 1.3080 ;
      RECT 2.0720 0.4200 2.3450 0.4700 ;
      RECT 2.1030 1.3080 2.3050 1.3580 ;
      RECT 2.2550 0.3710 2.3050 0.4200 ;
      RECT 2.1030 1.1660 2.1530 1.3080 ;
      RECT 2.8240 0.6040 3.4610 0.6540 ;
      RECT 2.8240 0.6540 2.8740 0.9780 ;
      RECT 2.5190 0.9780 2.8740 1.0270 ;
      RECT 2.5420 1.0270 2.8740 1.0280 ;
      RECT 2.5190 0.5880 2.5690 0.9780 ;
      RECT 2.8240 1.0280 2.8740 1.0290 ;
      RECT 2.5190 0.5380 2.6490 0.5880 ;
      RECT 2.7700 1.5210 3.1570 1.5710 ;
      RECT 1.4190 1.4780 1.7890 1.5280 ;
      RECT 1.4190 1.5280 1.4690 1.5650 ;
      RECT 1.0850 0.0960 1.4910 0.1460 ;
      RECT 1.2670 1.4280 1.3170 1.5260 ;
      RECT 1.2670 1.3780 1.9250 1.4280 ;
      RECT 1.8750 1.4280 1.9250 1.5840 ;
      RECT 0.7850 1.5260 1.3170 1.5760 ;
      RECT 0.5830 0.6180 1.0290 0.6680 ;
      RECT 0.5830 0.6680 0.6330 0.9140 ;
      RECT 0.5830 0.4220 0.6330 0.6180 ;
      RECT 1.0390 0.5180 1.1650 0.5680 ;
      RECT 1.0390 0.3940 1.0890 0.5180 ;
      RECT 1.1150 0.5680 1.1650 0.7180 ;
      RECT 1.0390 0.7180 1.1650 0.7680 ;
      RECT 1.0390 0.7680 1.0890 0.9140 ;
      RECT 2.9340 0.7090 3.1570 0.7590 ;
      RECT 2.5310 1.1490 2.5810 1.2720 ;
      RECT 2.3550 1.2720 2.5810 1.3220 ;
      RECT 2.3550 1.3220 2.4050 1.5220 ;
      RECT 2.1630 1.5220 2.4050 1.5720 ;
      RECT 2.9340 0.7590 2.9840 1.0990 ;
      RECT 2.5310 1.0990 2.9840 1.1490 ;
    LAYER PO ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 2.3410 0.7900 2.3710 1.6060 ;
      RECT 3.1010 0.0680 3.1310 0.7870 ;
      RECT 1.2770 0.0680 1.3070 0.5420 ;
      RECT 1.7330 0.0680 1.7630 0.6180 ;
      RECT 2.3410 0.0680 2.3710 0.6220 ;
      RECT 1.2770 0.7900 1.3070 1.6060 ;
      RECT 3.1010 1.0120 3.1310 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 1.7330 0.7300 1.7630 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 3.7090 0.0680 3.7390 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
  END
END DFFNX1_LVT

MACRO DFFNX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.256 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4710 0.1480 3.5210 0.3940 ;
        RECT 3.4710 0.3940 4.0170 0.4440 ;
        RECT 3.8970 0.4440 4.0170 0.5110 ;
        RECT 3.9670 0.5110 4.0170 0.8040 ;
        RECT 3.4710 0.8040 4.0170 0.8540 ;
        RECT 3.4710 0.8540 3.5210 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0490 0.0970 4.1590 0.2070 ;
        RECT 4.0910 0.2070 4.1410 0.2700 ;
        RECT 3.7750 0.2700 4.1410 0.3200 ;
        RECT 3.7750 0.1480 3.8250 0.2700 ;
        RECT 4.0910 0.3200 4.1410 0.9180 ;
        RECT 3.7750 0.9180 4.1410 0.9680 ;
        RECT 3.7750 0.9680 3.8250 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.2560 0.0300 ;
        RECT 0.5860 0.0300 0.6360 0.1960 ;
        RECT 1.7990 0.0300 1.8490 0.1990 ;
        RECT 3.9270 0.0300 3.9770 0.2200 ;
        RECT 3.6230 0.0300 3.6730 0.3190 ;
        RECT 3.3190 0.0300 3.3690 0.4080 ;
        RECT 0.2790 0.0300 0.3290 0.4190 ;
        RECT 3.1670 0.0300 3.2170 0.3300 ;
        RECT 0.5860 0.1960 0.9370 0.2460 ;
        RECT 1.7990 0.1990 2.0240 0.2490 ;
        RECT 2.6950 0.3300 3.2330 0.3800 ;
        RECT 0.8870 0.2460 0.9370 0.4500 ;
        RECT 0.7350 0.2460 0.7850 0.4500 ;
        RECT 1.7990 0.2490 1.8490 0.3730 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.2560 1.7020 ;
        RECT 0.2790 1.0330 0.3290 1.6420 ;
        RECT 3.3190 0.9120 3.3690 1.6420 ;
        RECT 3.6230 0.9600 3.6730 1.6420 ;
        RECT 3.9270 1.0520 3.9770 1.6420 ;
        RECT 2.6390 1.3580 2.6890 1.6420 ;
        RECT 1.9750 1.3280 2.0250 1.6420 ;
        RECT 3.2070 1.3580 3.2570 1.6420 ;
        RECT 0.4330 1.3540 0.4830 1.6420 ;
        RECT 2.6390 1.3080 2.7770 1.3580 ;
        RECT 1.7820 1.2780 2.0250 1.3280 ;
        RECT 3.1490 1.3080 3.2570 1.3580 ;
        RECT 0.4330 1.3340 0.9370 1.3540 ;
        RECT 0.4340 1.3040 0.9370 1.3340 ;
        RECT 0.7350 1.0880 0.7850 1.3040 ;
        RECT 0.8870 1.1010 0.9370 1.3040 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.3590 0.6800 ;
        RECT 0.2490 0.6800 0.4210 0.7300 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.4240 0.7250 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 4.3710 1.7730 ;
    LAYER M1 ;
      RECT 1.1910 0.2990 1.2810 0.3810 ;
      RECT 1.2150 0.3810 1.2650 0.9880 ;
      RECT 1.1910 1.0380 1.2410 1.3140 ;
      RECT 0.4310 0.9880 1.2650 1.0380 ;
      RECT 0.4310 1.0380 0.4810 1.2160 ;
      RECT 0.4310 0.8290 0.4810 0.9880 ;
      RECT 0.4310 0.5790 0.5210 0.6290 ;
      RECT 0.4310 0.4550 0.4810 0.5790 ;
      RECT 0.4310 0.7800 0.5210 0.8290 ;
      RECT 0.4710 0.6290 0.5210 0.7800 ;
      RECT 2.7870 0.1470 2.8370 0.2300 ;
      RECT 2.1150 0.2300 2.8370 0.2800 ;
      RECT 2.3150 0.1780 2.3970 0.2300 ;
      RECT 2.1150 0.2800 2.1650 0.3140 ;
      RECT 1.9640 0.3140 2.1650 0.3640 ;
      RECT 1.9640 0.3640 2.0140 0.5400 ;
      RECT 1.7070 0.5400 2.0140 0.5900 ;
      RECT 1.3430 0.6400 2.0930 0.6900 ;
      RECT 1.3430 0.6900 1.3930 1.1580 ;
      RECT 1.3430 0.4840 1.3930 0.6400 ;
      RECT 1.3430 1.1580 1.5610 1.2080 ;
      RECT 1.3430 0.4340 1.5610 0.4840 ;
      RECT 1.3430 1.2080 1.3930 1.3140 ;
      RECT 1.3430 0.3550 1.3930 0.4340 ;
      RECT 3.6800 0.6040 3.9170 0.6540 ;
      RECT 3.2070 0.7540 3.2570 1.2080 ;
      RECT 2.7100 0.5460 2.7600 0.6990 ;
      RECT 2.7100 0.4880 2.7600 0.4960 ;
      RECT 2.8470 1.2080 3.2570 1.2580 ;
      RECT 2.6190 0.6990 2.7600 0.7490 ;
      RECT 2.4070 0.4380 2.7600 0.4880 ;
      RECT 2.4070 0.4880 2.4570 1.1650 ;
      RECT 3.6800 0.6540 3.7300 0.7040 ;
      RECT 3.6800 0.5460 3.7300 0.6040 ;
      RECT 2.7100 0.4960 3.7300 0.5460 ;
      RECT 3.2070 0.7040 3.7300 0.7540 ;
      RECT 3.6800 0.4940 3.7300 0.4960 ;
      RECT 1.7070 0.7580 2.2290 0.8080 ;
      RECT 2.1790 0.5870 2.2290 0.7580 ;
      RECT 1.5500 1.0010 2.3450 1.0510 ;
      RECT 2.2950 0.4700 2.3450 1.0010 ;
      RECT 2.2550 1.0510 2.3050 1.3080 ;
      RECT 2.0720 0.4200 2.3450 0.4700 ;
      RECT 2.1030 1.3080 2.3050 1.3580 ;
      RECT 2.2550 0.3710 2.3050 0.4200 ;
      RECT 2.1030 1.1660 2.1530 1.3080 ;
      RECT 2.8240 0.6040 3.6130 0.6540 ;
      RECT 2.8240 0.6540 2.8740 0.9780 ;
      RECT 2.5190 0.9780 2.8740 1.0270 ;
      RECT 2.5420 1.0270 2.8740 1.0280 ;
      RECT 2.5190 0.5880 2.5690 0.9780 ;
      RECT 2.8240 1.0280 2.8740 1.0290 ;
      RECT 2.5190 0.5380 2.6490 0.5880 ;
      RECT 2.7700 1.5210 3.1570 1.5710 ;
      RECT 1.4190 1.4780 1.7890 1.5280 ;
      RECT 1.4190 1.5280 1.4690 1.5650 ;
      RECT 1.0850 0.0960 1.4910 0.1460 ;
      RECT 1.2670 1.4280 1.3170 1.5260 ;
      RECT 1.2670 1.3780 1.9250 1.4280 ;
      RECT 1.8750 1.4280 1.9250 1.5580 ;
      RECT 0.7850 1.5260 1.3170 1.5760 ;
      RECT 0.5830 0.6180 1.0290 0.6680 ;
      RECT 0.5830 0.6680 0.6330 0.9140 ;
      RECT 0.5830 0.4220 0.6330 0.6180 ;
      RECT 1.0390 0.5180 1.1650 0.5680 ;
      RECT 1.0390 0.3940 1.0890 0.5180 ;
      RECT 1.1150 0.5680 1.1650 0.7180 ;
      RECT 1.0390 0.7180 1.1650 0.7680 ;
      RECT 1.0390 0.7680 1.0890 0.9140 ;
      RECT 2.9340 0.7090 3.1570 0.7590 ;
      RECT 2.5310 1.1490 2.5810 1.2720 ;
      RECT 2.3550 1.2720 2.5810 1.3220 ;
      RECT 2.3550 1.3220 2.4050 1.5220 ;
      RECT 2.1630 1.5220 2.4050 1.5720 ;
      RECT 2.9340 0.7590 2.9840 1.0990 ;
      RECT 2.5310 1.0990 2.9840 1.1490 ;
    LAYER PO ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 1.7330 0.7300 1.7630 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 2.3410 0.7900 2.3710 1.6060 ;
      RECT 3.1010 0.0680 3.1310 0.7870 ;
      RECT 1.2770 0.0680 1.3070 0.5420 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 1.7330 0.0680 1.7630 0.6180 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 2.3410 0.0680 2.3710 0.6220 ;
      RECT 1.2770 0.7900 1.3070 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 3.7090 0.0680 3.7390 1.6060 ;
      RECT 3.1010 1.0120 3.1310 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
  END
END DFFNX2_LVT

MACRO DFFSSRX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.408 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.4080 1.7020 ;
        RECT 3.9270 0.9470 3.9770 1.6420 ;
        RECT 1.4050 1.3660 1.4550 1.6420 ;
        RECT 0.2790 1.3460 0.3290 1.6420 ;
        RECT 2.4070 1.3660 2.4570 1.6420 ;
        RECT 3.6630 1.4660 3.7130 1.6420 ;
        RECT 1.3050 1.3160 1.4550 1.3660 ;
        RECT 0.2790 1.2960 0.6330 1.3460 ;
        RECT 2.2550 1.3160 2.4570 1.3660 ;
        RECT 3.1510 1.4160 3.7130 1.4660 ;
        RECT 0.2790 0.9300 0.3290 1.2960 ;
        RECT 0.5830 0.9800 0.6330 1.2960 ;
        RECT 2.2550 1.1000 2.3050 1.3160 ;
        RECT 3.6230 1.1920 3.6730 1.4160 ;
    END
  END VDD

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0490 0.4270 4.1590 0.5110 ;
        RECT 3.7750 0.3770 4.1590 0.4270 ;
        RECT 4.1090 0.5110 4.1590 0.8080 ;
        RECT 3.7750 0.1360 3.8250 0.3770 ;
        RECT 3.7750 0.8080 4.1590 0.8580 ;
        RECT 3.7750 0.8580 3.8250 1.5460 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0790 1.0690 4.3110 1.1190 ;
        RECT 4.2010 1.0090 4.3110 1.0690 ;
        RECT 4.0790 1.1190 4.1290 1.5460 ;
        RECT 4.2610 0.3100 4.3110 1.0090 ;
        RECT 4.0790 0.2600 4.3110 0.3100 ;
        RECT 4.0790 0.1360 4.1290 0.2600 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7010 0.4210 0.7510 ;
        RECT 0.2490 0.7510 0.3590 0.8250 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END SETB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.4650 1.3330 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.4080 0.0300 ;
        RECT 3.1270 0.0300 3.1770 0.2040 ;
        RECT 0.2790 0.0300 0.3290 0.3550 ;
        RECT 3.9270 0.0300 3.9770 0.3030 ;
        RECT 3.6230 0.0300 3.6730 0.4010 ;
        RECT 2.0270 0.0300 2.0770 0.3010 ;
        RECT 3.1270 0.2040 3.2330 0.2540 ;
        RECT 0.2790 0.3550 0.6330 0.4050 ;
        RECT 1.3430 0.3010 2.4570 0.3510 ;
        RECT 0.5830 0.4050 0.6330 0.5290 ;
        RECT 0.2790 0.4050 0.3290 0.5130 ;
        RECT 2.4070 0.3510 2.4570 0.4750 ;
        RECT 1.3430 0.3510 1.3930 0.5760 ;
        RECT 2.2550 0.3510 2.3050 0.4750 ;
    END
  END VSS

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9470 0.8670 1.1190 0.9770 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 0.2010 0.7250 0.2510 ;
        RECT 0.4010 0.1070 0.5110 0.2010 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END RSTB
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 4.5230 1.7730 ;
    LAYER M1 ;
      RECT 1.0990 0.1040 1.9410 0.1540 ;
      RECT 1.7230 0.1540 1.7730 0.2170 ;
      RECT 1.0990 0.6260 1.4850 0.6760 ;
      RECT 1.1910 0.6760 1.2410 1.1520 ;
      RECT 1.1910 0.4010 1.2410 0.6260 ;
      RECT 1.8590 1.4170 2.2450 1.4670 ;
      RECT 0.4910 1.4490 0.8770 1.4990 ;
      RECT 1.4950 0.7260 1.5970 0.7760 ;
      RECT 1.4950 0.7760 1.5450 1.1520 ;
      RECT 1.5470 0.6760 1.5970 0.7260 ;
      RECT 1.5470 0.6260 1.6370 0.6760 ;
      RECT 1.5470 0.4960 1.5970 0.6260 ;
      RECT 1.4790 0.4460 1.5970 0.4960 ;
      RECT 3.8510 0.5270 3.9010 0.6580 ;
      RECT 3.2790 0.4770 3.9010 0.5270 ;
      RECT 2.8630 0.3000 2.9130 1.2160 ;
      RECT 3.2790 0.5270 3.3290 0.6540 ;
      RECT 3.0750 0.6540 3.3290 0.6770 ;
      RECT 3.0750 0.6770 3.4090 0.7040 ;
      RECT 3.2790 0.7040 3.4090 0.7270 ;
      RECT 3.3590 0.7270 3.4090 1.2160 ;
      RECT 2.8630 1.2160 3.4090 1.2660 ;
      RECT 1.6470 0.7260 1.7370 0.7760 ;
      RECT 1.6870 0.5760 1.7370 0.7260 ;
      RECT 1.6470 0.7760 1.6970 1.2020 ;
      RECT 1.6470 0.5260 1.7370 0.5760 ;
      RECT 0.8870 1.2020 1.6970 1.2520 ;
      RECT 1.6470 0.4300 1.6970 0.5260 ;
      RECT 0.8870 1.0970 0.9370 1.2020 ;
      RECT 0.8470 1.0470 0.9370 1.0970 ;
      RECT 0.8470 0.7520 1.0060 0.8020 ;
      RECT 0.9560 0.4930 1.0060 0.7520 ;
      RECT 0.8710 0.4430 1.0060 0.4930 ;
      RECT 0.8470 0.8020 0.8970 1.0470 ;
      RECT 2.8570 0.1040 3.0050 0.1510 ;
      RECT 2.1630 0.1510 3.0050 0.1540 ;
      RECT 2.1630 0.1540 2.9070 0.2010 ;
      RECT 0.7000 0.5730 0.8770 0.6230 ;
      RECT 0.7000 0.6230 0.7500 0.8440 ;
      RECT 0.4310 0.8440 0.7500 0.8940 ;
      RECT 0.4310 0.8940 0.4810 1.2460 ;
      RECT 0.4310 0.4550 0.4810 0.6010 ;
      RECT 0.4710 0.6510 0.5210 0.8440 ;
      RECT 0.4310 0.6010 0.5210 0.6510 ;
      RECT 2.0060 0.7730 2.7610 0.8230 ;
      RECT 2.7110 0.8230 2.7610 1.3800 ;
      RECT 2.5590 0.8230 2.6090 1.1660 ;
      RECT 2.7110 0.5020 2.7610 0.7730 ;
      RECT 2.5590 0.4520 2.7610 0.5020 ;
      RECT 2.5590 0.3000 2.6090 0.4520 ;
      RECT 2.7110 0.3000 2.7610 0.4520 ;
      RECT 3.5230 0.6770 3.6130 0.7270 ;
      RECT 3.5230 0.7270 3.5730 1.3160 ;
      RECT 2.8110 1.3160 3.5730 1.3660 ;
      RECT 2.8110 1.3660 2.8610 1.5280 ;
      RECT 2.5670 1.5280 2.8610 1.5780 ;
      RECT 2.5670 1.2660 2.6170 1.5280 ;
      RECT 2.4030 1.0440 2.4530 1.2160 ;
      RECT 2.1630 0.9940 2.4530 1.0440 ;
      RECT 2.4030 1.2160 2.6170 1.2660 ;
      RECT 1.7990 0.5730 2.5490 0.6230 ;
      RECT 1.9510 0.4300 2.0010 0.5730 ;
      RECT 1.7990 0.6230 1.8490 1.1960 ;
      RECT 1.7990 0.4300 1.8490 0.5730 ;
      RECT 1.7990 1.1960 2.0010 1.2460 ;
      RECT 1.9510 1.0720 2.0010 1.1960 ;
      RECT 3.7510 0.7080 4.0530 0.7580 ;
      RECT 4.0030 0.6210 4.0530 0.7080 ;
      RECT 3.7510 0.6270 3.8010 0.7080 ;
      RECT 3.3790 0.5770 3.8010 0.6270 ;
      RECT 2.9230 1.5280 3.6130 1.5780 ;
      RECT 3.3280 0.1540 3.3780 0.3040 ;
      RECT 2.9750 0.3040 3.3780 0.3540 ;
      RECT 3.2270 0.1040 3.4610 0.1540 ;
      RECT 2.9750 0.3540 3.0250 0.8080 ;
      RECT 2.9750 0.8080 3.0650 0.8580 ;
      RECT 3.0150 0.8580 3.0650 1.1660 ;
      RECT 0.7190 0.3010 1.1050 0.3510 ;
      RECT 0.7350 1.3160 1.1060 1.3660 ;
      RECT 0.7350 0.9800 0.7850 1.3160 ;
      RECT 1.8990 0.6730 2.2450 0.7230 ;
      RECT 1.8990 0.8800 2.1010 0.9300 ;
      RECT 2.0510 0.9300 2.1010 1.3170 ;
      RECT 1.8990 0.7230 1.9490 0.8800 ;
      RECT 1.7590 1.3170 2.1010 1.3670 ;
      RECT 1.7590 1.3670 1.8090 1.5280 ;
      RECT 1.5550 1.5280 1.8090 1.5780 ;
    LAYER PO ;
      RECT 3.7090 0.0760 3.7390 1.6060 ;
      RECT 0.8210 0.0760 0.8510 0.6510 ;
      RECT 1.7330 0.9200 1.7630 1.6060 ;
      RECT 1.5810 0.0760 1.6110 1.6060 ;
      RECT 2.0370 0.0760 2.0670 1.6060 ;
      RECT 3.8610 0.0760 3.8910 1.6060 ;
      RECT 1.4290 0.0760 1.4590 1.6060 ;
      RECT 2.4930 0.0760 2.5230 1.6060 ;
      RECT 0.0610 0.0760 0.0910 1.6060 ;
      RECT 3.5570 1.1320 3.5870 1.6060 ;
      RECT 2.1890 0.0760 2.2190 0.7510 ;
      RECT 3.1010 0.0760 3.1310 1.6060 ;
      RECT 3.4050 0.0760 3.4350 1.6060 ;
      RECT 1.8850 0.0760 1.9150 1.6060 ;
      RECT 4.0130 0.0760 4.0430 1.6060 ;
      RECT 3.2530 0.0760 3.2830 1.6060 ;
      RECT 1.1250 0.0760 1.1550 1.6060 ;
      RECT 2.7970 0.0760 2.8270 0.5970 ;
      RECT 2.6450 0.0760 2.6750 1.6060 ;
      RECT 0.6690 0.0760 0.6990 0.5970 ;
      RECT 0.6690 0.8160 0.6990 1.6060 ;
      RECT 2.9490 0.0760 2.9790 1.6060 ;
      RECT 0.9730 0.0760 1.0030 1.6060 ;
      RECT 0.2130 0.0760 0.2430 1.6060 ;
      RECT 0.3650 0.0760 0.3950 1.6060 ;
      RECT 2.1890 0.9660 2.2190 1.6060 ;
      RECT 1.2770 0.0760 1.3070 1.6060 ;
      RECT 4.3170 0.0760 4.3470 1.6060 ;
      RECT 2.3410 0.0760 2.3710 1.6060 ;
      RECT 0.8210 0.8700 0.8510 1.6060 ;
      RECT 1.7330 0.0760 1.7630 0.5970 ;
      RECT 2.7970 1.0320 2.8270 1.6060 ;
      RECT 4.1650 0.0760 4.1950 1.6060 ;
      RECT 0.5170 0.0760 0.5470 1.6060 ;
      RECT 3.5570 0.0760 3.5870 0.7550 ;
  END
END DFFSSRX1_LVT

MACRO CLOAD1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.76 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 0.7600 1.7020 ;
        RECT 0.4310 0.8230 0.4810 1.6420 ;
        RECT 0.2790 0.9150 0.3290 1.6420 ;
    END
  END VDD

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6600 0.4360 0.7100 ;
        RECT 0.2490 0.7100 0.3590 0.8150 ;
    END
  END A

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 0.7600 0.0300 ;
        RECT 0.4310 0.0300 0.4810 0.5020 ;
        RECT 0.2790 0.0300 0.3290 0.5020 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 0.8750 1.7730 ;
    LAYER PO ;
      RECT 0.3650 0.0690 0.3950 1.6060 ;
      RECT 0.2130 0.0710 0.2430 1.6060 ;
      RECT 0.6690 0.0710 0.6990 1.6060 ;
      RECT 0.5170 0.0710 0.5470 1.6060 ;
      RECT 0.0610 0.0710 0.0910 1.6060 ;
  END
END CLOAD1_LVT

MACRO DCAP_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.76 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 0.7600 1.7020 ;
        RECT 0.2790 1.2830 0.3290 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 0.7600 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.4870 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 0.8750 1.7730 ;
    LAYER M1 ;
      RECT 0.2350 1.1710 0.4810 1.2210 ;
      RECT 0.4310 1.2210 0.4810 1.5490 ;
      RECT 0.2350 0.6370 0.2850 1.1710 ;
      RECT 0.2350 0.5870 0.4360 0.6370 ;
      RECT 0.3390 1.0600 0.6210 1.1100 ;
      RECT 0.5710 0.3790 0.6210 1.0600 ;
      RECT 0.4310 0.3290 0.6210 0.3790 ;
      RECT 0.4310 0.3790 0.4810 0.4870 ;
      RECT 0.4310 0.1290 0.4810 0.3290 ;
    LAYER PO ;
      RECT 0.2130 0.0710 0.2430 1.6060 ;
      RECT 0.6690 0.0710 0.6990 1.6060 ;
      RECT 0.5170 0.0710 0.5470 1.6060 ;
      RECT 0.0610 0.0710 0.0910 1.6060 ;
      RECT 0.3650 0.0690 0.3950 0.6410 ;
      RECT 0.3650 1.0370 0.3950 1.6060 ;
  END
END DCAP_LVT

MACRO DEC24X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.648 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7070 1.4180 2.5320 1.4680 ;
        RECT 2.0730 1.4680 2.1830 1.5750 ;
        RECT 2.4820 1.4680 2.5320 1.5340 ;
        RECT 2.4820 1.5340 2.8530 1.5840 ;
    END
    ANTENNAGATEAREA 0.0732 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6430 1.5310 1.9530 1.5810 ;
        RECT 1.3320 1.4650 1.5190 1.5310 ;
    END
    ANTENNAGATEAREA 0.0732 ;
  END A1

  PIN Y2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2980 0.7650 3.4140 0.8150 ;
        RECT 3.3640 0.6630 3.4140 0.7650 ;
        RECT 3.3640 0.5530 3.5700 0.6630 ;
        RECT 3.3640 0.5450 3.4140 0.5530 ;
        RECT 3.2980 0.4950 3.4140 0.5450 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y2

  PIN Y3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1160 0.9900 0.3030 1.1320 ;
        RECT 0.2390 0.8300 0.2890 0.9900 ;
        RECT 0.2390 0.7800 0.3500 0.8300 ;
        RECT 0.2390 0.5410 0.2890 0.7800 ;
        RECT 0.2390 0.4910 0.3500 0.5410 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y3

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.6480 1.7020 ;
        RECT 3.1670 1.3470 3.2170 1.6420 ;
        RECT 0.4310 1.3350 0.4810 1.6420 ;
        RECT 2.6950 1.2970 3.2330 1.3470 ;
        RECT 0.4090 1.2850 2.4800 1.3350 ;
    END
  END VDD

  PIN Y0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0630 0.8350 2.1750 0.8850 ;
        RECT 2.0630 0.5450 2.1130 0.8350 ;
        RECT 2.0630 0.5110 2.1970 0.5450 ;
        RECT 2.0630 0.4950 2.2870 0.5110 ;
        RECT 2.0920 0.4010 2.2870 0.4950 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y0

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.6480 0.0300 ;
        RECT 3.1670 0.0300 3.2170 0.1370 ;
        RECT 0.4310 0.0300 0.4810 0.1370 ;
        RECT 0.4310 0.1370 3.2400 0.1460 ;
        RECT 1.3490 0.0960 1.8890 0.1370 ;
        RECT 0.4310 0.1460 1.4130 0.1870 ;
        RECT 1.8390 0.1460 3.2400 0.1870 ;
        RECT 0.4310 0.1870 0.4810 0.2160 ;
        RECT 1.8390 0.1870 1.8890 0.3570 ;
        RECT 1.7800 0.3570 1.8890 0.4070 ;
    END
  END VSS

  PIN Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3320 0.8570 1.5690 0.9670 ;
        RECT 1.5190 0.5410 1.5690 0.8570 ;
        RECT 1.4740 0.4910 1.5690 0.5410 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y1
  OBS
    LAYER NWELL ;
      RECT -0.0700 0.6790 3.7180 1.7730 ;
    LAYER M1 ;
      RECT 2.5820 1.4310 2.7010 1.4810 ;
      RECT 2.5820 1.2350 2.6320 1.4310 ;
      RECT 0.8880 1.1850 2.6320 1.2350 ;
      RECT 1.6190 0.4600 1.6970 0.5420 ;
      RECT 1.6190 0.5420 1.6690 1.1850 ;
      RECT 0.8880 0.8380 0.9380 1.1850 ;
      RECT 0.8880 0.7880 1.0320 0.8380 ;
      RECT 1.1910 0.6520 1.4690 0.7020 ;
      RECT 1.4190 0.7020 1.4690 0.7220 ;
      RECT 1.4190 0.6240 1.4690 0.6520 ;
      RECT 1.1910 0.4600 1.2410 0.6520 ;
      RECT 1.1910 0.7020 1.2410 0.9810 ;
      RECT 1.0190 0.9810 1.2410 1.0310 ;
      RECT 1.5760 0.1960 1.7890 0.2460 ;
      RECT 1.5760 0.2460 1.6260 0.3600 ;
      RECT 0.8110 0.3600 1.6260 0.4100 ;
      RECT 0.8110 0.4100 0.8610 0.6610 ;
      RECT 2.3410 0.9810 2.6250 1.0310 ;
      RECT 2.3410 0.7050 2.3910 0.9810 ;
      RECT 2.1630 0.6550 2.3910 0.7050 ;
      RECT 2.3410 0.5260 2.3910 0.6550 ;
      RECT 2.3410 0.4760 2.4730 0.5260 ;
      RECT 2.4830 0.8810 2.7250 0.9310 ;
      RECT 2.6750 0.9310 2.7250 1.0810 ;
      RECT 2.4830 0.6680 2.5330 0.8810 ;
      RECT 1.9510 1.0810 2.7250 1.1310 ;
      RECT 2.4830 0.6180 3.0050 0.6680 ;
      RECT 2.4830 0.6020 2.5340 0.6180 ;
      RECT 1.9510 0.4600 2.0010 1.0810 ;
      RECT 3.0550 0.6510 3.3140 0.7010 ;
      RECT 3.0550 0.7010 3.1050 1.0100 ;
      RECT 3.0550 0.5260 3.1050 0.6510 ;
      RECT 2.8470 1.0100 3.1050 1.0600 ;
      RECT 2.9940 0.4760 3.1050 0.5260 ;
      RECT 0.5830 0.9810 0.8010 1.0310 ;
      RECT 0.5830 0.7050 0.6330 0.9810 ;
      RECT 0.3390 0.6550 0.6330 0.7050 ;
      RECT 0.5830 0.4600 0.6330 0.6550 ;
    LAYER PO ;
      RECT 1.1250 0.0670 1.1550 1.6090 ;
      RECT 0.2130 0.0700 0.2430 1.6090 ;
      RECT 1.7330 0.0710 1.7630 1.6090 ;
      RECT 2.7970 0.0710 2.8270 1.6090 ;
      RECT 3.1010 0.0710 3.1310 1.6090 ;
      RECT 0.5170 0.0710 0.5470 1.6090 ;
      RECT 0.0610 0.0700 0.0910 1.6090 ;
      RECT 0.9730 0.0710 1.0030 1.6090 ;
      RECT 2.6450 0.0710 2.6750 1.6090 ;
      RECT 2.1890 0.0710 2.2190 1.6090 ;
      RECT 2.0370 0.0710 2.0670 1.6090 ;
      RECT 2.4930 0.0710 2.5230 1.6090 ;
      RECT 0.6690 0.0710 0.6990 1.6090 ;
      RECT 0.8210 0.0710 0.8510 1.6090 ;
      RECT 1.2770 0.0710 1.3070 1.6090 ;
      RECT 1.8850 0.0710 1.9150 1.6090 ;
      RECT 3.4050 0.0710 3.4350 1.6090 ;
      RECT 2.3410 0.0710 2.3710 1.6090 ;
      RECT 3.5570 0.0710 3.5870 1.6090 ;
      RECT 1.5810 0.0710 1.6110 1.6090 ;
      RECT 2.9490 0.0710 2.9790 1.6090 ;
      RECT 3.2530 0.0710 3.2830 1.6090 ;
      RECT 0.3650 0.0710 0.3950 1.6090 ;
      RECT 1.4290 0.0710 1.4590 1.6090 ;
  END
END DEC24X1_LVT

MACRO DEC24X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.256 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0110 1.4180 2.9880 1.4680 ;
        RECT 2.3770 1.4680 2.4870 1.5750 ;
        RECT 2.9380 1.4680 2.9880 1.5340 ;
        RECT 2.9380 1.5340 3.3090 1.5840 ;
    END
    ANTENNAGATEAREA 0.0732 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7890 1.5310 2.2570 1.5810 ;
        RECT 1.7330 1.4650 1.8780 1.5310 ;
    END
    ANTENNAGATEAREA 0.0732 ;
  END A1

  PIN Y2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.7540 0.7650 4.0850 0.8150 ;
        RECT 4.0350 0.6630 4.0850 0.7650 ;
        RECT 4.0350 0.5530 4.1780 0.6630 ;
        RECT 4.0350 0.5450 4.0850 0.5530 ;
        RECT 3.7540 0.4950 4.0850 0.5450 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Y2

  PIN Y3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2390 0.8300 0.2890 0.9900 ;
        RECT 0.2390 0.9900 0.3780 1.1320 ;
        RECT 0.2390 0.7800 0.5020 0.8300 ;
        RECT 0.2390 0.5410 0.2890 0.7800 ;
        RECT 0.2390 0.4910 0.5020 0.5410 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Y3

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.2560 1.7020 ;
        RECT 3.6230 1.3470 3.6730 1.6420 ;
        RECT 0.5830 1.3350 0.6330 1.6420 ;
        RECT 3.1510 1.2970 3.9930 1.3470 ;
        RECT 0.2630 1.2860 2.9290 1.3350 ;
        RECT 1.5210 1.3350 2.9290 1.3360 ;
        RECT 0.2630 1.2850 1.5650 1.2860 ;
    END
  END VDD

  PIN Y0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3670 0.8350 2.6310 0.8850 ;
        RECT 2.3670 0.5450 2.4170 0.8350 ;
        RECT 2.3670 0.5110 2.6300 0.5450 ;
        RECT 2.3670 0.4950 2.6580 0.5110 ;
        RECT 2.5290 0.4010 2.6580 0.4950 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Y0

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.2560 0.0300 ;
        RECT 3.6230 0.0300 3.6730 0.1370 ;
        RECT 0.5830 0.0300 0.6330 0.1370 ;
        RECT 0.2630 0.1370 3.9930 0.1460 ;
        RECT 1.8010 0.0960 2.1930 0.1370 ;
        RECT 0.2630 0.1460 1.8650 0.1870 ;
        RECT 2.1430 0.1460 3.9930 0.1870 ;
        RECT 0.5830 0.1870 0.6330 0.2160 ;
        RECT 2.1430 0.1870 2.1930 0.3570 ;
        RECT 2.0840 0.3570 2.1930 0.4070 ;
    END
  END VSS

  PIN Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6170 0.8570 1.8730 0.9670 ;
        RECT 1.8230 0.5410 1.8730 0.8570 ;
        RECT 1.6260 0.4910 1.8730 0.5410 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Y1
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 4.3710 1.7730 ;
    LAYER M1 ;
      RECT 3.0380 1.4340 3.1570 1.4840 ;
      RECT 3.0380 1.2350 3.0880 1.4340 ;
      RECT 1.0400 1.1850 3.0880 1.2350 ;
      RECT 1.9230 0.4600 2.0010 0.5420 ;
      RECT 1.9230 0.5420 1.9730 1.1850 ;
      RECT 1.0400 0.8380 1.0900 1.1850 ;
      RECT 1.0400 0.7880 1.1840 0.8380 ;
      RECT 1.3430 0.6520 1.7730 0.7020 ;
      RECT 1.7230 0.7020 1.7730 0.7220 ;
      RECT 1.7230 0.6240 1.7730 0.6520 ;
      RECT 1.5710 0.7020 1.6210 0.7220 ;
      RECT 1.5710 0.6240 1.6210 0.6520 ;
      RECT 1.3430 0.7020 1.3930 0.9810 ;
      RECT 1.3430 0.4600 1.3930 0.6520 ;
      RECT 1.1710 0.9810 1.3930 1.0310 ;
      RECT 1.9160 0.1960 2.0930 0.2460 ;
      RECT 1.9160 0.2460 1.9660 0.3600 ;
      RECT 0.9630 0.3600 1.9660 0.4100 ;
      RECT 0.9630 0.4100 1.0130 0.6610 ;
      RECT 2.7970 0.9810 3.0810 1.0310 ;
      RECT 2.7970 0.6890 2.8470 0.9810 ;
      RECT 2.4670 0.6390 2.8470 0.6890 ;
      RECT 2.7970 0.5260 2.8470 0.6390 ;
      RECT 2.7970 0.4760 2.9290 0.5260 ;
      RECT 2.9390 0.8810 3.1810 0.9310 ;
      RECT 3.1310 0.9310 3.1810 1.0810 ;
      RECT 2.9390 0.6680 2.9890 0.8810 ;
      RECT 2.2550 1.0810 3.1810 1.1310 ;
      RECT 2.9390 0.6180 3.4610 0.6680 ;
      RECT 2.9390 0.6020 2.9900 0.6180 ;
      RECT 2.2550 0.4600 2.3050 1.0810 ;
      RECT 3.5110 0.6260 3.9170 0.6760 ;
      RECT 3.5110 0.6760 3.5610 1.0100 ;
      RECT 3.5110 0.5260 3.5610 0.6260 ;
      RECT 3.3030 1.0100 3.5610 1.0600 ;
      RECT 3.4500 0.4760 3.5610 0.5260 ;
      RECT 0.7350 0.9810 0.9530 1.0310 ;
      RECT 0.7350 0.6970 0.7850 0.9810 ;
      RECT 0.3390 0.6470 0.7850 0.6970 ;
      RECT 0.7350 0.4600 0.7850 0.6470 ;
    LAYER PO ;
      RECT 1.8850 0.0710 1.9150 1.6090 ;
      RECT 3.2530 0.0710 3.2830 1.6090 ;
      RECT 3.5570 0.0710 3.5870 1.6090 ;
      RECT 0.6690 0.0710 0.6990 1.6090 ;
      RECT 1.7330 0.0710 1.7630 1.6090 ;
      RECT 1.4290 0.0670 1.4590 1.6090 ;
      RECT 0.3650 0.0710 0.3950 1.6090 ;
      RECT 0.5170 0.0700 0.5470 1.6090 ;
      RECT 2.0370 0.0710 2.0670 1.6090 ;
      RECT 3.1010 0.0710 3.1310 1.6090 ;
      RECT 3.4050 0.0710 3.4350 1.6090 ;
      RECT 0.8210 0.0710 0.8510 1.6090 ;
      RECT 1.2770 0.0710 1.3070 1.6090 ;
      RECT 2.9490 0.0710 2.9790 1.6090 ;
      RECT 2.4930 0.0710 2.5230 1.6090 ;
      RECT 2.3410 0.0710 2.3710 1.6090 ;
      RECT 0.0610 0.0710 0.0910 1.6090 ;
      RECT 0.2130 0.0710 0.2430 1.6090 ;
      RECT 4.0130 0.0710 4.0430 1.6090 ;
      RECT 4.1650 0.0710 4.1950 1.6090 ;
      RECT 2.7970 0.0710 2.8270 1.6090 ;
      RECT 0.9730 0.0710 1.0030 1.6090 ;
      RECT 1.1250 0.0710 1.1550 1.6090 ;
      RECT 1.5810 0.0710 1.6110 1.6090 ;
      RECT 2.1890 0.0710 2.2190 1.6090 ;
      RECT 3.7090 0.0710 3.7390 1.6090 ;
      RECT 2.6450 0.0710 2.6750 1.6090 ;
      RECT 3.8610 0.0710 3.8910 1.6090 ;
  END
END DEC24X2_LVT

MACRO DELLN1X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.04 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0970 0.6750 0.4210 0.7250 ;
        RECT 0.0970 0.7250 0.2100 0.8150 ;
    END
    ANTENNAGATEAREA 0.0105 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.0400 1.7020 ;
        RECT 1.4950 1.1500 1.5450 1.6420 ;
        RECT 0.5830 1.2900 0.6330 1.6420 ;
        RECT 1.1910 0.7970 1.2410 1.6420 ;
        RECT 2.1030 0.8160 2.1530 1.6420 ;
        RECT 0.2790 0.8170 0.3290 1.6420 ;
        RECT 2.5590 0.9920 2.6090 1.6420 ;
        RECT 1.4550 1.1000 1.5450 1.1500 ;
        RECT 0.5430 1.2400 0.6330 1.2900 ;
        RECT 1.4550 0.9500 1.5050 1.1000 ;
        RECT 0.5430 1.0900 0.5930 1.2400 ;
        RECT 1.4550 0.9000 1.5490 0.9500 ;
        RECT 0.5430 1.0400 0.6210 1.0900 ;
        RECT 1.4990 0.6490 1.5490 0.9000 ;
        RECT 0.5710 0.6190 0.6210 1.0400 ;
        RECT 1.4990 0.5990 1.7890 0.6490 ;
        RECT 0.5710 0.5690 0.8770 0.6190 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.0400 0.0300 ;
        RECT 1.9910 0.0300 2.0410 0.1980 ;
        RECT 1.0790 0.0300 1.1290 0.1980 ;
        RECT 2.1030 0.0300 2.1530 0.5470 ;
        RECT 0.2790 0.0300 0.3290 0.5400 ;
        RECT 2.5590 0.0300 2.6090 0.4100 ;
        RECT 1.1910 0.0300 1.2410 0.5500 ;
        RECT 1.4950 0.1980 2.0410 0.2480 ;
        RECT 0.5830 0.1980 1.1290 0.2480 ;
        RECT 1.4950 0.2480 1.5450 0.4990 ;
        RECT 0.5830 0.2480 0.6330 0.4690 ;
        RECT 1.4950 0.4990 1.8890 0.5490 ;
        RECT 0.5830 0.4690 0.9770 0.5190 ;
        RECT 1.8390 0.5490 1.8890 1.0000 ;
        RECT 0.9270 0.5190 0.9770 1.1400 ;
        RECT 1.5550 1.0000 1.8890 1.0500 ;
        RECT 0.6430 1.1400 0.9770 1.1900 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4070 0.1310 2.4570 0.5370 ;
        RECT 2.4070 0.5370 2.9430 0.5870 ;
        RECT 2.7510 0.5870 2.9430 0.6630 ;
        RECT 2.7110 0.1310 2.7610 0.5370 ;
        RECT 2.7510 0.6630 2.8010 0.8920 ;
        RECT 2.4070 0.8920 2.8010 0.9420 ;
        RECT 2.7110 0.9420 2.7610 1.5490 ;
        RECT 2.4070 0.9420 2.4570 1.5490 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 3.1650 1.7730 ;
    LAYER M1 ;
      RECT 1.0390 0.6750 1.3330 0.7250 ;
      RECT 1.0390 0.7250 1.0890 1.5340 ;
      RECT 1.0390 0.3470 1.0890 0.6750 ;
      RECT 0.4310 0.0960 1.0290 0.1460 ;
      RECT 0.4310 0.7750 0.5210 0.8250 ;
      RECT 0.4310 0.5410 0.5210 0.5910 ;
      RECT 0.4710 0.5910 0.5210 0.7750 ;
      RECT 0.4310 0.1460 0.4810 0.5410 ;
      RECT 0.4310 0.8250 0.4810 0.9990 ;
      RECT 1.9510 0.6600 2.2450 0.7100 ;
      RECT 1.9510 0.7100 2.0010 1.5370 ;
      RECT 1.9510 0.3710 2.0010 0.6600 ;
      RECT 1.3430 0.0960 1.9410 0.1460 ;
      RECT 1.3430 0.1460 1.3930 0.5320 ;
      RECT 1.3430 0.8250 1.3930 0.9710 ;
      RECT 1.3430 0.5320 1.4330 0.5820 ;
      RECT 1.3830 0.5820 1.4330 0.7750 ;
      RECT 1.3430 0.7750 1.4330 0.8250 ;
      RECT 2.2950 0.6600 2.7010 0.7100 ;
      RECT 2.2950 0.7100 2.3450 0.8870 ;
      RECT 2.2950 0.5820 2.3450 0.6600 ;
      RECT 2.2550 0.8870 2.3450 0.9370 ;
      RECT 2.2550 0.5320 2.3450 0.5820 ;
      RECT 2.2550 0.9370 2.3050 1.2690 ;
      RECT 2.2550 0.2810 2.3050 0.5320 ;
    LAYER PO ;
      RECT 1.7330 0.0660 1.7630 0.6830 ;
      RECT 1.5810 0.0660 1.6110 0.6830 ;
      RECT 1.5810 0.9700 1.6110 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.6690 1.1100 0.6990 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 2.4930 0.0660 2.5230 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 2.6450 0.0660 2.6750 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 0.8210 0.0660 0.8510 0.6530 ;
      RECT 0.6690 0.0660 0.6990 0.6530 ;
      RECT 0.8210 1.1100 0.8510 1.6060 ;
      RECT 1.7330 0.9700 1.7630 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
  END
END DELLN1X2_LVT

MACRO DELLN2X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.952 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0970 0.6750 0.4210 0.7250 ;
        RECT 0.0970 0.7250 0.2100 0.8150 ;
    END
    ANTENNAGATEAREA 0.0102 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.9520 1.7020 ;
        RECT 3.4710 0.9920 3.5210 1.6420 ;
        RECT 2.1030 0.7750 2.1530 1.6420 ;
        RECT 0.5830 1.2100 0.6330 1.6420 ;
        RECT 1.4950 1.2900 1.5450 1.6420 ;
        RECT 1.1910 0.8170 1.2410 1.6420 ;
        RECT 3.0150 0.8160 3.0650 1.6420 ;
        RECT 0.2790 0.8070 0.3290 1.6420 ;
        RECT 2.3670 1.4280 2.4170 1.6420 ;
        RECT 0.5430 1.1600 0.6330 1.2100 ;
        RECT 1.4550 1.2400 1.5450 1.2900 ;
        RECT 2.3670 1.3780 2.4570 1.4280 ;
        RECT 0.5430 1.0100 0.5930 1.1600 ;
        RECT 1.4550 1.0910 1.5050 1.2400 ;
        RECT 2.4070 0.6490 2.4570 1.3780 ;
        RECT 0.5430 0.9600 0.6370 1.0100 ;
        RECT 1.4550 1.0410 1.5450 1.0910 ;
        RECT 2.4070 0.5990 2.7010 0.6490 ;
        RECT 0.5870 0.6490 0.6370 0.9600 ;
        RECT 1.4950 0.6490 1.5450 1.0410 ;
        RECT 0.5870 0.5990 0.8770 0.6490 ;
        RECT 1.4950 0.5990 1.7890 0.6490 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.3190 0.5370 3.8550 0.5870 ;
        RECT 3.3190 0.1160 3.3690 0.5370 ;
        RECT 3.6790 0.5870 3.8550 0.6630 ;
        RECT 3.6230 0.1160 3.6730 0.5370 ;
        RECT 3.6790 0.6630 3.7290 0.8920 ;
        RECT 3.3190 0.8920 3.7290 0.9420 ;
        RECT 3.6230 0.9420 3.6730 1.5640 ;
        RECT 3.3190 0.9420 3.3690 1.5640 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END Y

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.9520 0.0300 ;
        RECT 1.9910 0.0300 2.0410 0.1980 ;
        RECT 3.4710 0.0300 3.5210 0.4100 ;
        RECT 2.1060 0.0300 2.1560 0.2660 ;
        RECT 2.9030 0.0300 2.9530 0.1980 ;
        RECT 1.0790 0.0300 1.1290 0.1980 ;
        RECT 1.1910 0.0300 1.2410 0.5400 ;
        RECT 3.0150 0.0300 3.0650 0.5470 ;
        RECT 0.2790 0.0300 0.3290 0.5400 ;
        RECT 1.4950 0.1980 2.0410 0.2480 ;
        RECT 2.1030 0.2660 2.1560 0.3160 ;
        RECT 2.4070 0.1980 2.9530 0.2480 ;
        RECT 0.5830 0.1980 1.1290 0.2480 ;
        RECT 1.4950 0.2480 1.5450 0.4990 ;
        RECT 2.1030 0.3160 2.1530 0.5800 ;
        RECT 2.4070 0.2480 2.4570 0.4990 ;
        RECT 0.5830 0.2480 0.6330 0.4990 ;
        RECT 1.4950 0.4990 1.8890 0.5490 ;
        RECT 2.4070 0.4990 2.8010 0.5490 ;
        RECT 0.5830 0.4990 0.9770 0.5490 ;
        RECT 1.8390 0.5490 1.8890 1.1400 ;
        RECT 2.7510 0.5490 2.8010 1.5220 ;
        RECT 0.9270 0.5490 0.9770 1.0600 ;
        RECT 1.5550 1.1400 1.8890 1.1900 ;
        RECT 2.4670 1.5220 2.8010 1.5720 ;
        RECT 0.6430 1.0600 0.9770 1.1100 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 4.0670 1.7730 ;
    LAYER M1 ;
      RECT 3.2070 0.6600 3.6280 0.7100 ;
      RECT 3.2070 0.7100 3.2570 0.8870 ;
      RECT 3.2070 0.5820 3.2570 0.6600 ;
      RECT 3.1670 0.8870 3.2570 0.9370 ;
      RECT 3.1670 0.5320 3.2570 0.5820 ;
      RECT 3.1670 0.9370 3.2170 1.2660 ;
      RECT 3.1670 0.2850 3.2170 0.5320 ;
      RECT 2.8630 0.6600 3.1570 0.7100 ;
      RECT 2.8630 0.7100 2.9130 1.4300 ;
      RECT 2.8630 0.3770 2.9130 0.6600 ;
      RECT 2.2550 0.0960 2.8530 0.1460 ;
      RECT 2.2550 0.1460 2.3050 0.5320 ;
      RECT 2.2550 0.5320 2.3450 0.5820 ;
      RECT 2.2950 0.5820 2.3450 0.7750 ;
      RECT 2.2550 0.7750 2.3450 0.8250 ;
      RECT 2.2550 0.8250 2.3050 0.8870 ;
      RECT 1.0390 0.6750 1.3330 0.7250 ;
      RECT 1.0390 0.7250 1.0890 1.5050 ;
      RECT 1.0390 0.3770 1.0890 0.6750 ;
      RECT 0.4310 0.0960 1.0290 0.1460 ;
      RECT 0.4310 0.1460 0.4810 0.5410 ;
      RECT 0.4310 0.8250 0.4810 0.9640 ;
      RECT 0.4310 0.5410 0.5210 0.5910 ;
      RECT 0.4710 0.5910 0.5210 0.7750 ;
      RECT 0.4310 0.7750 0.5210 0.8250 ;
      RECT 1.9510 0.6710 2.2450 0.7210 ;
      RECT 1.9510 0.7210 2.0010 1.4930 ;
      RECT 1.9510 0.3810 2.0010 0.6710 ;
      RECT 1.3430 0.0960 1.9410 0.1460 ;
      RECT 1.3430 0.1460 1.3930 0.5320 ;
      RECT 1.3430 0.5320 1.4330 0.5820 ;
      RECT 1.3830 0.5820 1.4330 0.7750 ;
      RECT 1.3430 0.7750 1.4330 0.8250 ;
      RECT 1.3430 0.8250 1.3930 0.9910 ;
    LAYER PO ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 2.4930 0.0660 2.5230 0.6830 ;
      RECT 2.4930 0.8260 2.5230 1.6060 ;
      RECT 2.6450 0.0660 2.6750 0.6830 ;
      RECT 2.6450 0.8260 2.6750 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 0.8210 0.0660 0.8510 0.6830 ;
      RECT 0.6690 0.0660 0.6990 0.6830 ;
      RECT 0.8210 1.0300 0.8510 1.6060 ;
      RECT 1.7330 1.1100 1.7630 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 1.7330 0.0660 1.7630 0.6830 ;
      RECT 1.5810 0.0660 1.6110 0.6830 ;
      RECT 1.5810 1.1100 1.6110 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 3.5570 0.0660 3.5870 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 3.7090 0.0660 3.7390 1.6060 ;
      RECT 3.4050 0.0660 3.4350 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 0.6690 1.0300 0.6990 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
  END
END DELLN2X2_LVT

MACRO DELLN3X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.776 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0970 0.6750 0.4210 0.7250 ;
        RECT 0.0970 0.7250 0.2100 0.8150 ;
    END
    ANTENNAGATEAREA 0.0096 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 5.7760 1.7020 ;
        RECT 4.1910 1.4280 4.2410 1.6420 ;
        RECT 4.1910 1.3780 4.2810 1.4280 ;
        RECT 2.4070 1.3300 2.4570 1.6420 ;
        RECT 2.3670 1.2800 2.4570 1.3300 ;
        RECT 3.3190 1.2700 3.3690 1.6420 ;
        RECT 3.2790 1.2200 3.3690 1.2700 ;
        RECT 0.5830 1.2100 0.6330 1.6420 ;
        RECT 1.4950 1.2100 1.5450 1.6420 ;
        RECT 1.4550 1.1600 1.5450 1.2100 ;
        RECT 0.5430 1.1600 0.6330 1.2100 ;
        RECT 2.3670 1.1300 2.4170 1.2800 ;
        RECT 2.3670 1.0800 2.4610 1.1300 ;
        RECT 3.2790 1.0710 3.3290 1.2200 ;
        RECT 3.2790 1.0210 3.3690 1.0710 ;
        RECT 5.2950 0.9920 5.3450 1.6420 ;
        RECT 1.4550 1.0100 1.5050 1.1600 ;
        RECT 0.5430 0.9890 0.5930 1.1600 ;
        RECT 1.4550 0.9600 1.5490 1.0100 ;
        RECT 3.0150 0.8170 3.0650 1.6420 ;
        RECT 3.9270 0.7750 3.9770 1.6420 ;
        RECT 4.8390 0.8160 4.8890 1.6420 ;
        RECT 4.2310 0.6490 4.2810 1.3780 ;
        RECT 3.3190 0.6490 3.3690 1.0210 ;
        RECT 4.2310 0.5990 4.5250 0.6490 ;
        RECT 3.3190 0.5990 3.6130 0.6490 ;
        RECT 1.1910 0.7950 1.2410 1.6420 ;
        RECT 0.2790 0.7950 0.3290 1.6420 ;
        RECT 2.1030 0.8070 2.1530 1.6420 ;
        RECT 2.4110 0.6490 2.4610 1.0800 ;
        RECT 0.5430 0.9390 0.6370 0.9890 ;
        RECT 1.4990 0.6490 1.5490 0.9600 ;
        RECT 0.5870 0.6490 0.6370 0.9390 ;
        RECT 2.4110 0.5990 2.7010 0.6490 ;
        RECT 1.4990 0.5990 1.7890 0.6490 ;
        RECT 0.5870 0.5990 0.8770 0.6490 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.1430 0.5370 5.6790 0.5870 ;
        RECT 5.1430 0.1160 5.1930 0.5370 ;
        RECT 5.5030 0.5870 5.6790 0.6630 ;
        RECT 5.4470 0.1160 5.4970 0.5370 ;
        RECT 5.5030 0.6630 5.5530 0.8920 ;
        RECT 5.1430 0.8920 5.5530 0.9420 ;
        RECT 5.4470 0.9420 5.4970 1.5640 ;
        RECT 5.1430 0.9420 5.1930 1.5640 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END Y

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 4.2910 1.5220 4.6250 1.5720 ;
        RECT 2.4670 1.1800 2.8010 1.2300 ;
        RECT 3.3790 1.1200 3.7130 1.1700 ;
        RECT 1.5550 1.0600 1.8890 1.1100 ;
        RECT 0.6430 1.0400 0.9770 1.0900 ;
        RECT 4.5750 0.5490 4.6250 1.5220 ;
        RECT 2.7510 0.5490 2.8010 1.1800 ;
        RECT 3.6630 0.5490 3.7130 1.1200 ;
        RECT 1.8390 0.5490 1.8890 1.0600 ;
        RECT 0.9270 0.5490 0.9770 1.0400 ;
        RECT 4.2310 0.4990 4.6250 0.5490 ;
        RECT 3.3190 0.4990 3.7130 0.5490 ;
        RECT 0.5830 0.4990 0.9770 0.5490 ;
        RECT 1.4950 0.4990 1.8890 0.5490 ;
        RECT 2.4070 0.4990 2.8010 0.5490 ;
        RECT 3.9270 0.3160 3.9770 0.5800 ;
        RECT 3.9270 0.2660 3.9800 0.3160 ;
        RECT 4.2310 0.2480 4.2810 0.4990 ;
        RECT 3.3190 0.2480 3.3690 0.4990 ;
        RECT 0.5830 0.2480 0.6330 0.4990 ;
        RECT 1.4950 0.2480 1.5450 0.4990 ;
        RECT 2.4070 0.2480 2.4570 0.4990 ;
        RECT 2.4070 0.1980 2.9530 0.2480 ;
        RECT 0.0000 -0.0300 5.7760 0.0300 ;
        RECT 4.8390 0.0300 4.8890 0.5470 ;
        RECT 3.0150 0.0300 3.0650 0.5400 ;
        RECT 5.2950 0.0300 5.3450 0.4100 ;
        RECT 3.9300 0.0300 3.9800 0.2660 ;
        RECT 4.2310 0.1980 4.7770 0.2480 ;
        RECT 3.3190 0.1980 3.8650 0.2480 ;
        RECT 3.8150 0.0300 3.8650 0.1980 ;
        RECT 2.9030 0.0300 2.9530 0.1980 ;
        RECT 4.7270 0.0300 4.7770 0.1980 ;
        RECT 0.2790 0.0300 0.3290 0.5600 ;
        RECT 1.1910 0.0300 1.2410 0.5600 ;
        RECT 2.1030 0.0300 2.1530 0.5400 ;
        RECT 0.5830 0.1980 1.1290 0.2480 ;
        RECT 1.4950 0.1980 2.0410 0.2480 ;
        RECT 1.9910 0.0300 2.0410 0.1980 ;
        RECT 1.0790 0.0300 1.1290 0.1980 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 5.8910 1.7730 ;
    LAYER M1 ;
      RECT 2.8630 0.6750 3.1570 0.7250 ;
      RECT 2.8630 0.7250 2.9130 1.5050 ;
      RECT 2.8630 0.3770 2.9130 0.6750 ;
      RECT 1.0390 0.6750 1.3330 0.7250 ;
      RECT 1.0390 0.7250 1.0890 1.5050 ;
      RECT 1.0390 0.3310 1.0890 0.6750 ;
      RECT 0.4310 0.0960 1.0290 0.1460 ;
      RECT 0.4310 0.1460 0.4810 0.5410 ;
      RECT 0.4310 0.5410 0.5210 0.5910 ;
      RECT 0.4310 0.8250 0.4810 0.8870 ;
      RECT 0.4710 0.5910 0.5210 0.7750 ;
      RECT 0.4310 0.7750 0.5210 0.8250 ;
      RECT 3.1670 0.0960 3.7650 0.1460 ;
      RECT 3.1670 0.1460 3.2170 0.5320 ;
      RECT 3.1670 0.5320 3.2570 0.5820 ;
      RECT 3.2070 0.5820 3.2570 0.7750 ;
      RECT 3.1670 0.7750 3.2570 0.8250 ;
      RECT 3.1670 0.8250 3.2170 0.9210 ;
      RECT 2.2550 0.0960 2.8530 0.1460 ;
      RECT 2.2550 0.1460 2.3050 0.5410 ;
      RECT 2.2550 0.5410 2.3450 0.5910 ;
      RECT 2.2950 0.5910 2.3450 0.7750 ;
      RECT 2.2550 0.7750 2.3450 0.8250 ;
      RECT 2.2550 0.8250 2.3050 0.8720 ;
      RECT 1.9510 0.6750 2.2450 0.7250 ;
      RECT 1.9510 0.7250 2.0010 1.5050 ;
      RECT 1.9510 0.3010 2.0010 0.6750 ;
      RECT 5.0310 0.6600 5.4520 0.7100 ;
      RECT 5.0310 0.7100 5.0810 0.8870 ;
      RECT 5.0310 0.5820 5.0810 0.6600 ;
      RECT 4.9910 0.8870 5.0810 0.9370 ;
      RECT 4.9910 0.5320 5.0810 0.5820 ;
      RECT 4.9910 0.9370 5.0410 1.2660 ;
      RECT 4.9910 0.2850 5.0410 0.5320 ;
      RECT 3.7750 0.6710 4.0690 0.7210 ;
      RECT 3.7750 0.7210 3.8250 1.4930 ;
      RECT 3.7750 0.3810 3.8250 0.6710 ;
      RECT 1.3430 0.0960 1.9410 0.1460 ;
      RECT 1.3430 0.1460 1.3930 0.5410 ;
      RECT 1.3430 0.5410 1.4330 0.5910 ;
      RECT 1.3830 0.5910 1.4330 0.7750 ;
      RECT 1.3430 0.7750 1.4330 0.8250 ;
      RECT 1.3430 0.8250 1.3930 0.8870 ;
      RECT 4.6870 0.6600 4.9810 0.7100 ;
      RECT 4.6870 0.7100 4.7370 1.4300 ;
      RECT 4.6870 0.3770 4.7370 0.6600 ;
      RECT 4.0790 0.0960 4.6770 0.1460 ;
      RECT 4.0790 0.1460 4.1290 0.5320 ;
      RECT 4.0790 0.5320 4.1690 0.5820 ;
      RECT 4.1190 0.5820 4.1690 0.7750 ;
      RECT 4.0790 0.7750 4.1690 0.8250 ;
      RECT 4.0790 0.8250 4.1290 0.8870 ;
    LAYER PO ;
      RECT 2.9490 0.0660 2.9790 1.6060 ;
      RECT 2.6450 0.0660 2.6750 0.6830 ;
      RECT 2.4930 0.0660 2.5230 0.6830 ;
      RECT 2.6450 1.1500 2.6750 1.6060 ;
      RECT 3.5570 1.0900 3.5870 1.6060 ;
      RECT 3.2530 0.0660 3.2830 1.6060 ;
      RECT 3.5570 0.0660 3.5870 0.6830 ;
      RECT 3.4050 0.0660 3.4350 0.6830 ;
      RECT 3.4050 1.0900 3.4350 1.6060 ;
      RECT 3.7090 0.0660 3.7390 1.6060 ;
      RECT 5.0770 0.0660 5.1070 1.6060 ;
      RECT 3.1010 0.0660 3.1310 1.6060 ;
      RECT 5.3810 0.0660 5.4110 1.6060 ;
      RECT 4.9250 0.0660 4.9550 1.6060 ;
      RECT 5.5330 0.0660 5.5630 1.6060 ;
      RECT 5.2290 0.0660 5.2590 1.6060 ;
      RECT 5.6850 0.0660 5.7150 1.6060 ;
      RECT 2.4930 1.1500 2.5230 1.6060 ;
      RECT 4.0130 0.0660 4.0430 1.6060 ;
      RECT 3.8610 0.0660 3.8910 1.6060 ;
      RECT 4.1650 0.0660 4.1950 1.6060 ;
      RECT 4.7730 0.0660 4.8030 1.6060 ;
      RECT 4.6210 0.0660 4.6510 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 0.6690 0.0660 0.6990 0.6830 ;
      RECT 0.8210 0.0660 0.8510 0.6830 ;
      RECT 0.6690 1.0100 0.6990 1.6060 ;
      RECT 0.8210 1.0100 0.8510 1.6060 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 1.8850 0.0660 1.9150 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 2.0370 0.0660 2.0670 1.6060 ;
      RECT 1.7330 0.0660 1.7630 0.6830 ;
      RECT 1.5810 0.0660 1.6110 0.6830 ;
      RECT 1.7330 1.0300 1.7630 1.6060 ;
      RECT 1.5810 1.0300 1.6110 1.6060 ;
      RECT 4.3170 0.0660 4.3470 0.6830 ;
      RECT 4.3170 0.9760 4.3470 1.6060 ;
      RECT 4.4690 0.0660 4.4990 0.6830 ;
      RECT 4.4690 0.9760 4.4990 1.6060 ;
      RECT 2.3410 0.0660 2.3710 1.6060 ;
      RECT 2.7970 0.0660 2.8270 1.6060 ;
      RECT 2.1890 0.0660 2.2190 1.6060 ;
  END
END DELLN3X2_LVT

MACRO DFFARX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.256 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.2560 0.0300 ;
        RECT 0.5860 0.0300 0.6360 0.1960 ;
        RECT 0.2790 0.0300 0.3290 0.4190 ;
        RECT 3.7750 0.0300 3.8250 0.2200 ;
        RECT 3.4710 0.0300 3.5210 0.3300 ;
        RECT 1.5410 0.0300 1.5910 0.2870 ;
        RECT 0.5860 0.1960 0.9370 0.2460 ;
        RECT 2.9990 0.3300 3.5370 0.3800 ;
        RECT 1.5410 0.2870 2.0010 0.3370 ;
        RECT 0.8870 0.2460 0.9370 0.4500 ;
        RECT 0.7350 0.2460 0.7850 0.4500 ;
        RECT 1.9510 0.3370 2.0010 0.4610 ;
        RECT 1.9510 0.2490 2.0010 0.2870 ;
        RECT 1.9510 0.1990 2.1760 0.2490 ;
    END
  END VSS

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0500 1.1610 4.1600 1.2210 ;
        RECT 3.9270 1.2210 4.1600 1.2710 ;
        RECT 4.1090 0.2040 4.1590 1.1610 ;
        RECT 3.9270 1.2710 3.9770 1.5460 ;
        RECT 3.9110 0.1540 4.1590 0.2040 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.2560 1.7020 ;
        RECT 0.2790 1.0330 0.3290 1.6420 ;
        RECT 3.7750 0.9470 3.8250 1.6420 ;
        RECT 2.1270 1.3280 2.1770 1.6420 ;
        RECT 3.5110 1.3580 3.5610 1.6420 ;
        RECT 0.8870 1.3640 0.9370 1.6420 ;
        RECT 1.9340 1.2780 2.1770 1.3280 ;
        RECT 2.8340 1.3080 3.5610 1.3580 ;
        RECT 0.7350 1.3140 0.9370 1.3640 ;
        RECT 0.7350 1.0980 0.7850 1.3140 ;
        RECT 0.8870 1.1110 0.9370 1.3140 ;
    END
  END VDD

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7230 0.0880 2.8530 0.1380 ;
        RECT 2.7710 0.1380 2.8530 0.1740 ;
        RECT 1.7230 0.1380 1.8790 0.2070 ;
    END
    ANTENNAGATEAREA 0.0441 ;
  END RSTB

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.3590 0.6800 ;
        RECT 0.2490 0.6800 0.4210 0.7300 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.4240 0.7250 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8970 1.0090 4.0070 1.1190 ;
        RECT 3.9570 0.8540 4.0070 1.0090 ;
        RECT 3.6230 0.8040 4.0070 0.8540 ;
        RECT 3.6230 0.8540 3.6730 1.5460 ;
        RECT 3.9570 0.3590 4.0070 0.8040 ;
        RECT 3.6230 0.3090 4.0070 0.3590 ;
        RECT 3.6230 0.1480 3.6730 0.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 4.3710 1.7730 ;
    LAYER M1 ;
      RECT 1.1910 0.2990 1.2810 0.3810 ;
      RECT 1.2150 0.3810 1.2650 0.9880 ;
      RECT 0.4310 0.9880 1.2650 1.0380 ;
      RECT 1.1910 1.0380 1.2410 1.3140 ;
      RECT 0.4310 1.0380 0.4810 1.2160 ;
      RECT 0.4310 0.8290 0.4810 0.9880 ;
      RECT 0.4310 0.5790 0.5210 0.6290 ;
      RECT 0.4310 0.4550 0.4810 0.5790 ;
      RECT 0.4310 0.7800 0.5210 0.8290 ;
      RECT 0.4710 0.6290 0.5210 0.7800 ;
      RECT 3.0910 0.0990 3.1410 0.2300 ;
      RECT 2.2490 0.2300 3.1410 0.2800 ;
      RECT 2.4670 0.2800 2.5490 0.2900 ;
      RECT 2.2490 0.2800 2.2990 0.3140 ;
      RECT 2.0980 0.3140 2.2990 0.3640 ;
      RECT 2.0980 0.3640 2.1480 0.5400 ;
      RECT 1.8590 0.5400 2.1480 0.5900 ;
      RECT 2.4670 0.1880 2.5490 0.2300 ;
      RECT 1.3430 0.6400 2.2450 0.6900 ;
      RECT 1.3430 0.6900 1.3930 1.1580 ;
      RECT 1.3430 0.4840 1.3930 0.6400 ;
      RECT 1.3430 1.2080 1.3930 1.3140 ;
      RECT 1.3430 0.3550 1.3930 0.4340 ;
      RECT 1.3430 1.1580 1.7130 1.2080 ;
      RECT 1.3430 0.4340 1.5610 0.4840 ;
      RECT 2.5590 0.4380 3.9010 0.4880 ;
      RECT 3.8510 0.4880 3.9010 0.7040 ;
      RECT 3.5110 0.7040 3.9010 0.7540 ;
      RECT 2.5590 0.4880 2.6090 1.1650 ;
      RECT 2.8620 0.4880 2.9120 0.7660 ;
      RECT 2.8620 0.7660 3.0050 0.8160 ;
      RECT 3.5110 0.7540 3.5610 1.2080 ;
      RECT 3.1510 1.2080 3.5610 1.2580 ;
      RECT 1.8590 0.7860 2.3810 0.8360 ;
      RECT 2.3310 0.6210 2.3810 0.7860 ;
      RECT 3.0550 0.6040 3.7650 0.6540 ;
      RECT 3.0550 0.6540 3.1050 0.9780 ;
      RECT 2.6940 0.9780 3.1050 1.0280 ;
      RECT 2.6940 0.5880 2.7440 0.9780 ;
      RECT 2.6940 0.5380 2.8010 0.5880 ;
      RECT 2.2550 1.3080 2.4570 1.3580 ;
      RECT 2.2550 1.1010 2.3050 1.3080 ;
      RECT 2.4070 1.0510 2.4570 1.3080 ;
      RECT 1.5500 1.0010 2.4970 1.0510 ;
      RECT 2.4470 0.5690 2.4970 1.0010 ;
      RECT 2.4070 0.5190 2.4970 0.5690 ;
      RECT 2.4070 0.4700 2.4570 0.5190 ;
      RECT 2.2240 0.4200 2.4570 0.4700 ;
      RECT 2.4070 0.3810 2.4570 0.4200 ;
      RECT 1.4190 1.4780 1.9410 1.5280 ;
      RECT 1.4190 1.5280 1.4690 1.5650 ;
      RECT 1.0870 1.5260 1.3170 1.5760 ;
      RECT 1.2670 1.4280 1.3170 1.5260 ;
      RECT 1.2670 1.3780 2.0770 1.4280 ;
      RECT 2.0270 1.4280 2.0770 1.5840 ;
      RECT 0.5830 0.6180 1.0290 0.6680 ;
      RECT 0.5830 0.6680 0.6330 0.9140 ;
      RECT 0.5830 0.4220 0.6330 0.6180 ;
      RECT 1.0390 0.5180 1.1650 0.5680 ;
      RECT 1.0390 0.3940 1.0890 0.5180 ;
      RECT 1.1150 0.5680 1.1650 0.7180 ;
      RECT 1.0390 0.7180 1.1650 0.7680 ;
      RECT 1.0390 0.7680 1.0890 0.9140 ;
      RECT 3.0740 1.4290 3.4610 1.4790 ;
      RECT 3.2380 0.7090 3.4610 0.7590 ;
      RECT 3.2380 0.7590 3.2880 1.0990 ;
      RECT 2.6830 1.0990 3.2880 1.1490 ;
      RECT 2.6830 1.1490 2.7330 1.2720 ;
      RECT 2.5070 1.2720 2.7330 1.3220 ;
      RECT 2.5070 1.3220 2.5570 1.5280 ;
      RECT 2.3150 1.5280 2.5570 1.5780 ;
      RECT 1.4790 1.2780 1.8650 1.3280 ;
      RECT 0.7810 0.0960 1.4910 0.1460 ;
    LAYER PO ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 3.7090 0.0680 3.7390 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 1.2770 0.0680 1.3070 0.5420 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 1.2770 0.9900 1.3070 1.6060 ;
      RECT 3.4050 1.0120 3.4350 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 1.8850 0.0680 1.9150 0.6180 ;
      RECT 3.4050 0.0680 3.4350 0.7870 ;
      RECT 2.4930 0.8820 2.5230 1.6060 ;
      RECT 2.4930 0.0680 2.5230 0.6320 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 1.8850 0.7580 1.9150 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
  END
END DFFARX1_LVT

MACRO DFFARX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.56 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.7750 0.8040 4.3210 0.8540 ;
        RECT 3.7750 0.8540 3.8250 1.5460 ;
        RECT 4.2710 0.5110 4.3210 0.8040 ;
        RECT 4.2010 0.4440 4.3210 0.5110 ;
        RECT 3.7750 0.3940 4.3210 0.4440 ;
        RECT 3.7750 0.1480 3.8250 0.3940 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.3530 0.0970 4.4630 0.2070 ;
        RECT 4.3950 0.2070 4.4450 0.2700 ;
        RECT 4.0790 0.2700 4.4450 0.3200 ;
        RECT 4.0790 0.1480 4.1290 0.2700 ;
        RECT 4.3950 0.3200 4.4450 0.9180 ;
        RECT 4.0790 0.9180 4.4450 0.9680 ;
        RECT 4.0790 0.9680 4.1290 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.5600 0.0300 ;
        RECT 0.5860 0.0300 0.6360 0.1960 ;
        RECT 1.5590 0.0300 1.6090 0.2870 ;
        RECT 4.2310 0.0300 4.2810 0.2200 ;
        RECT 3.9270 0.0300 3.9770 0.3190 ;
        RECT 3.6230 0.0300 3.6730 0.4080 ;
        RECT 0.2790 0.0300 0.3290 0.4190 ;
        RECT 3.4710 0.0300 3.5210 0.3300 ;
        RECT 0.5860 0.1960 0.9370 0.2460 ;
        RECT 1.5590 0.2870 2.0010 0.3370 ;
        RECT 2.9990 0.3300 3.5370 0.3800 ;
        RECT 0.8870 0.2460 0.9370 0.4500 ;
        RECT 0.7350 0.2460 0.7850 0.4500 ;
        RECT 1.9510 0.3370 2.0010 0.4610 ;
        RECT 1.9510 0.2490 2.0010 0.2870 ;
        RECT 1.9510 0.1990 2.1760 0.2490 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.5600 1.7020 ;
        RECT 0.2790 1.0330 0.3290 1.6420 ;
        RECT 3.6230 0.9120 3.6730 1.6420 ;
        RECT 3.9270 0.9600 3.9770 1.6420 ;
        RECT 4.2310 1.0520 4.2810 1.6420 ;
        RECT 2.1370 1.3280 2.1870 1.6420 ;
        RECT 3.5110 1.3580 3.5610 1.6420 ;
        RECT 0.8870 1.3640 0.9370 1.6420 ;
        RECT 1.9340 1.2780 2.1870 1.3280 ;
        RECT 2.8340 1.3080 3.5610 1.3580 ;
        RECT 0.7350 1.3140 0.9370 1.3640 ;
        RECT 0.7350 1.0980 0.7850 1.3140 ;
        RECT 0.8870 1.1110 0.9370 1.3140 ;
    END
  END VDD

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7230 0.0880 2.8530 0.1380 ;
        RECT 2.7710 0.1380 2.8530 0.1740 ;
        RECT 1.7230 0.1380 1.8790 0.2070 ;
    END
    ANTENNAGATEAREA 0.0441 ;
  END RSTB

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.3590 0.6800 ;
        RECT 0.2490 0.6800 0.4210 0.7300 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.4240 0.7250 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 4.6750 1.7730 ;
    LAYER M1 ;
      RECT 1.1910 0.2990 1.2810 0.3810 ;
      RECT 1.2150 0.3810 1.2650 0.9880 ;
      RECT 0.4310 0.9880 1.2650 1.0380 ;
      RECT 1.1910 1.0380 1.2410 1.3140 ;
      RECT 0.4310 1.0380 0.4810 1.2160 ;
      RECT 0.4310 0.8290 0.4810 0.9880 ;
      RECT 0.4310 0.5790 0.5210 0.6290 ;
      RECT 0.4310 0.4550 0.4810 0.5790 ;
      RECT 0.4310 0.7800 0.5210 0.8290 ;
      RECT 0.4710 0.6290 0.5210 0.7800 ;
      RECT 3.0910 0.0880 3.1410 0.2300 ;
      RECT 2.2490 0.2300 3.1410 0.2800 ;
      RECT 2.4670 0.2800 2.5490 0.2900 ;
      RECT 2.2490 0.2800 2.2990 0.3140 ;
      RECT 2.0980 0.3140 2.2990 0.3640 ;
      RECT 2.0980 0.3640 2.1480 0.5400 ;
      RECT 1.8590 0.5400 2.1480 0.5900 ;
      RECT 2.4670 0.1880 2.5490 0.2300 ;
      RECT 1.3430 0.6400 2.2450 0.6900 ;
      RECT 1.3430 0.6900 1.3930 1.1580 ;
      RECT 1.3430 0.4840 1.3930 0.6400 ;
      RECT 1.3430 1.2080 1.3930 1.3140 ;
      RECT 1.3430 0.3550 1.3930 0.4340 ;
      RECT 1.3430 1.1580 1.7130 1.2080 ;
      RECT 1.3430 0.4340 1.5610 0.4840 ;
      RECT 3.9840 0.6040 4.2210 0.6540 ;
      RECT 2.8620 0.5540 2.9120 0.7660 ;
      RECT 2.8620 0.4880 2.9120 0.5040 ;
      RECT 3.5110 0.7540 3.5610 1.2080 ;
      RECT 2.8620 0.7660 3.0050 0.8160 ;
      RECT 2.5590 0.4380 2.9120 0.4880 ;
      RECT 3.1510 1.2080 3.5610 1.2580 ;
      RECT 2.5590 0.4880 2.6090 1.1650 ;
      RECT 3.9840 0.5540 4.0340 0.6040 ;
      RECT 3.9840 0.6540 4.0340 0.7040 ;
      RECT 2.8620 0.5040 4.0340 0.5540 ;
      RECT 3.9840 0.5030 4.0340 0.5040 ;
      RECT 3.5110 0.7040 4.0340 0.7540 ;
      RECT 1.8590 0.7860 2.3810 0.8360 ;
      RECT 2.3310 0.6210 2.3810 0.7860 ;
      RECT 0.7810 0.0960 1.4910 0.1460 ;
      RECT 3.0550 0.6040 3.9170 0.6540 ;
      RECT 3.0550 0.6540 3.1050 0.9780 ;
      RECT 2.6940 0.9780 3.1050 1.0280 ;
      RECT 2.6940 0.5880 2.7440 0.9780 ;
      RECT 2.6940 0.5380 2.8010 0.5880 ;
      RECT 2.2550 1.3080 2.4570 1.3580 ;
      RECT 2.2550 1.1010 2.3050 1.3080 ;
      RECT 2.4070 1.0510 2.4570 1.3080 ;
      RECT 1.5500 1.0010 2.4970 1.0510 ;
      RECT 2.4470 0.5590 2.4970 1.0010 ;
      RECT 2.4070 0.5090 2.4970 0.5590 ;
      RECT 2.4070 0.4700 2.4570 0.5090 ;
      RECT 2.2240 0.4200 2.4570 0.4700 ;
      RECT 2.4070 0.3710 2.4570 0.4200 ;
      RECT 1.4190 1.4780 1.9410 1.5280 ;
      RECT 1.4190 1.5280 1.4690 1.5650 ;
      RECT 1.0870 1.5260 1.3170 1.5760 ;
      RECT 1.2670 1.4280 1.3170 1.5260 ;
      RECT 1.2670 1.3780 2.0770 1.4280 ;
      RECT 2.0270 1.4280 2.0770 1.5840 ;
      RECT 0.5830 0.6180 1.0290 0.6680 ;
      RECT 0.5830 0.6680 0.6330 0.9140 ;
      RECT 0.5830 0.4220 0.6330 0.6180 ;
      RECT 1.0390 0.5180 1.1650 0.5680 ;
      RECT 1.0390 0.3940 1.0890 0.5180 ;
      RECT 1.1150 0.5680 1.1650 0.7180 ;
      RECT 1.0390 0.7180 1.1650 0.7680 ;
      RECT 1.0390 0.7680 1.0890 0.9140 ;
      RECT 3.0740 1.4290 3.4610 1.4790 ;
      RECT 3.2380 0.7090 3.4610 0.7590 ;
      RECT 3.2380 0.7590 3.2880 1.0990 ;
      RECT 2.6830 1.0990 3.2880 1.1490 ;
      RECT 2.6830 1.1490 2.7330 1.2720 ;
      RECT 2.5070 1.2720 2.7330 1.3220 ;
      RECT 2.5070 1.3220 2.5570 1.5280 ;
      RECT 2.3150 1.5280 2.5570 1.5780 ;
      RECT 1.4790 1.2780 1.8650 1.3280 ;
    LAYER PO ;
      RECT 2.4930 0.0680 2.5230 0.6330 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 1.8850 0.7580 1.9150 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 1.2770 0.0680 1.3070 0.5420 ;
      RECT 1.2770 0.9900 1.3070 1.6060 ;
      RECT 3.4050 1.0120 3.4350 1.6060 ;
      RECT 3.7090 0.0680 3.7390 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 4.4690 0.0680 4.4990 1.6060 ;
      RECT 1.8850 0.0680 1.9150 0.6180 ;
      RECT 3.4050 0.0680 3.4350 0.7870 ;
      RECT 2.4930 0.8820 2.5230 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 4.3170 0.0680 4.3470 1.6060 ;
  END
END DFFARX2_LVT

MACRO DFFASRX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.56 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.5600 0.0300 ;
        RECT 0.5860 0.0300 0.6360 0.1960 ;
        RECT 0.2790 0.0300 0.3290 0.4190 ;
        RECT 4.0790 0.0300 4.1290 0.2200 ;
        RECT 1.5410 0.0300 1.5910 0.2870 ;
        RECT 3.7750 0.0300 3.8250 0.3300 ;
        RECT 0.5860 0.1960 0.9370 0.2460 ;
        RECT 1.5410 0.2870 2.1530 0.3370 ;
        RECT 3.1510 0.3300 3.8410 0.3800 ;
        RECT 0.8870 0.2460 0.9370 0.4500 ;
        RECT 0.7350 0.2460 0.7850 0.4500 ;
        RECT 2.1030 0.3370 2.1530 0.4610 ;
        RECT 1.9510 0.3370 2.0010 0.4610 ;
    END
  END VSS

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.3540 1.1610 4.4640 1.2210 ;
        RECT 4.2310 1.2210 4.4640 1.2710 ;
        RECT 4.4130 0.2040 4.4630 1.1610 ;
        RECT 4.2310 1.2710 4.2810 1.5460 ;
        RECT 4.2150 0.1540 4.4630 0.2040 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.5600 1.7020 ;
        RECT 0.2790 1.0330 0.3290 1.6420 ;
        RECT 4.0790 0.9470 4.1290 1.6420 ;
        RECT 0.8870 1.3540 0.9370 1.6420 ;
        RECT 2.1270 1.3280 2.1770 1.6420 ;
        RECT 3.8150 1.3580 3.8650 1.6420 ;
        RECT 0.7350 1.3040 0.9370 1.3540 ;
        RECT 1.9340 1.2780 2.3360 1.3280 ;
        RECT 2.9860 1.3080 3.8650 1.3580 ;
        RECT 0.7350 1.0880 0.7850 1.3040 ;
        RECT 0.8870 1.1010 0.9370 1.3040 ;
    END
  END VDD

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9230 0.1430 3.0050 0.1790 ;
        RECT 1.7230 0.0930 3.0050 0.1430 ;
        RECT 1.7230 0.1430 1.8790 0.2070 ;
    END
    ANTENNAGATEAREA 0.0441 ;
  END RSTB

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.3590 0.6800 ;
        RECT 0.2490 0.6800 0.4210 0.7300 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.5310 0.8570 3.7030 1.0340 ;
    END
    ANTENNAGATEAREA 0.0441 ;
  END SETB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.4240 0.7250 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.2010 1.0090 4.3110 1.1190 ;
        RECT 4.2610 0.8540 4.3110 1.0090 ;
        RECT 3.9270 0.8040 4.3110 0.8540 ;
        RECT 3.9270 0.8540 3.9770 1.5460 ;
        RECT 4.2610 0.3590 4.3110 0.8040 ;
        RECT 3.9270 0.3090 4.3110 0.3590 ;
        RECT 3.9270 0.1480 3.9770 0.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 4.6750 1.7730 ;
    LAYER M1 ;
      RECT 1.1910 0.2990 1.2810 0.3810 ;
      RECT 1.2150 0.3810 1.2650 0.9880 ;
      RECT 1.1910 1.0380 1.2410 1.3140 ;
      RECT 0.4310 0.9880 1.2650 1.0380 ;
      RECT 0.4310 1.0380 0.4810 1.2160 ;
      RECT 0.4310 0.8290 0.4810 0.9880 ;
      RECT 0.4310 0.5790 0.5210 0.6290 ;
      RECT 0.4310 0.4550 0.4810 0.5790 ;
      RECT 0.4310 0.7800 0.5210 0.8290 ;
      RECT 0.4710 0.6290 0.5210 0.7800 ;
      RECT 3.2430 0.0880 3.2930 0.2300 ;
      RECT 2.2950 0.2300 3.2930 0.2800 ;
      RECT 2.6190 0.2800 2.7010 0.2950 ;
      RECT 2.2950 0.2800 2.3450 0.5400 ;
      RECT 1.8590 0.5400 2.3450 0.5900 ;
      RECT 2.6190 0.1930 2.7010 0.2300 ;
      RECT 1.3430 0.6400 2.2450 0.6900 ;
      RECT 1.3430 0.6900 1.3930 1.1580 ;
      RECT 1.3430 0.4840 1.3930 0.6400 ;
      RECT 1.3430 1.2080 1.3930 1.3140 ;
      RECT 1.3430 0.3550 1.3930 0.4340 ;
      RECT 1.3430 1.1580 1.7130 1.2080 ;
      RECT 1.3430 0.4340 1.5610 0.4840 ;
      RECT 1.8590 0.7860 2.5490 0.8360 ;
      RECT 4.1550 0.4880 4.2050 0.7040 ;
      RECT 2.7110 0.4380 4.2050 0.4880 ;
      RECT 3.8150 0.7040 4.2050 0.7540 ;
      RECT 3.8150 0.7540 3.8650 1.1080 ;
      RECT 3.4550 1.1080 3.8650 1.1580 ;
      RECT 2.7110 0.4880 2.7610 1.1650 ;
      RECT 3.0140 0.4880 3.0640 0.7660 ;
      RECT 3.0140 0.7660 3.1570 0.8160 ;
      RECT 2.5590 0.6210 2.6490 0.6710 ;
      RECT 2.5990 0.6710 2.6490 1.0010 ;
      RECT 2.5590 0.4960 2.6090 0.6210 ;
      RECT 1.5500 1.0010 2.6490 1.0510 ;
      RECT 2.4070 0.4460 2.6090 0.4960 ;
      RECT 2.5590 1.0510 2.6090 1.3080 ;
      RECT 2.4070 0.3710 2.4570 0.4460 ;
      RECT 2.5590 0.3860 2.6090 0.4460 ;
      RECT 2.4070 1.3080 2.6090 1.3580 ;
      RECT 2.4070 1.2160 2.4570 1.3080 ;
      RECT 2.0860 1.1660 2.4570 1.2160 ;
      RECT 3.2070 0.6040 4.0690 0.6540 ;
      RECT 3.2070 0.6540 3.2570 0.9780 ;
      RECT 2.8460 0.9780 3.2570 1.0280 ;
      RECT 2.8460 0.5880 2.8960 0.9780 ;
      RECT 2.8460 0.5380 2.9530 0.5880 ;
      RECT 3.2260 1.4080 3.7650 1.4580 ;
      RECT 1.4190 1.4780 1.9410 1.5280 ;
      RECT 1.4190 1.5280 1.4690 1.5650 ;
      RECT 1.0990 1.5260 1.3170 1.5760 ;
      RECT 1.2670 1.4280 1.3170 1.5260 ;
      RECT 1.2670 1.3780 2.0770 1.4280 ;
      RECT 2.0270 1.4280 2.0770 1.5440 ;
      RECT 0.5830 0.6180 1.0290 0.6680 ;
      RECT 0.5830 0.6680 0.6330 0.9140 ;
      RECT 0.5830 0.4220 0.6330 0.6180 ;
      RECT 1.0390 0.5180 1.1650 0.5680 ;
      RECT 1.0390 0.3940 1.0890 0.5180 ;
      RECT 1.1150 0.5680 1.1650 0.7180 ;
      RECT 1.0390 0.7180 1.1650 0.7680 ;
      RECT 1.0390 0.7680 1.0890 0.9140 ;
      RECT 3.3450 0.7090 3.7650 0.7590 ;
      RECT 3.3450 0.7590 3.3950 1.0990 ;
      RECT 2.8350 1.0990 3.3950 1.1490 ;
      RECT 2.8350 1.1490 2.8850 1.2720 ;
      RECT 2.6590 1.2720 2.8850 1.3220 ;
      RECT 2.6590 1.3220 2.7090 1.4280 ;
      RECT 2.4670 1.4280 2.7090 1.4780 ;
      RECT 0.7950 0.0960 1.4910 0.1460 ;
      RECT 2.2860 1.5280 3.6260 1.5780 ;
      RECT 3.3030 1.2080 3.6890 1.2580 ;
      RECT 1.4790 1.2780 1.8650 1.3280 ;
    LAYER PO ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 1.2770 0.0680 1.3070 0.5420 ;
      RECT 4.4690 0.0680 4.4990 1.6060 ;
      RECT 1.2770 0.9900 1.3070 1.6060 ;
      RECT 3.7090 0.0680 3.7390 0.7870 ;
      RECT 1.8850 0.0680 1.9150 0.6180 ;
      RECT 2.6450 0.8820 2.6750 1.6060 ;
      RECT 3.7090 1.0120 3.7390 1.6060 ;
      RECT 2.6450 0.0680 2.6750 0.6370 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 1.8850 0.7580 1.9150 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 4.3170 0.0680 4.3470 1.6060 ;
  END
END DFFASRX1_LVT

MACRO DFFASRX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.864 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0790 0.3940 4.5870 0.4010 ;
        RECT 4.0790 0.1480 4.1290 0.3940 ;
        RECT 4.0790 0.4010 4.6250 0.4440 ;
        RECT 4.5050 0.4440 4.6250 0.5110 ;
        RECT 4.5750 0.5110 4.6250 0.8040 ;
        RECT 4.0790 0.8040 4.6250 0.8540 ;
        RECT 4.5750 0.8540 4.6250 0.8610 ;
        RECT 4.0790 0.8540 4.1290 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.6570 0.2170 4.7670 0.2700 ;
        RECT 4.3830 0.2700 4.7670 0.3200 ;
        RECT 4.6570 0.3200 4.7670 0.3590 ;
        RECT 4.3830 0.1480 4.4330 0.2700 ;
        RECT 4.6990 0.3590 4.7490 0.9180 ;
        RECT 4.3830 0.9180 4.7490 0.9680 ;
        RECT 4.3830 0.9680 4.4330 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.8640 0.0300 ;
        RECT 0.5860 0.0300 0.6360 0.1960 ;
        RECT 4.5350 0.0300 4.5850 0.2200 ;
        RECT 4.2310 0.0300 4.2810 0.3190 ;
        RECT 3.9270 0.0300 3.9770 0.4080 ;
        RECT 0.2790 0.0300 0.3290 0.4190 ;
        RECT 1.5410 0.0300 1.5910 0.2870 ;
        RECT 3.7750 0.0300 3.8250 0.3300 ;
        RECT 0.5860 0.1960 0.9370 0.2460 ;
        RECT 1.5410 0.2870 2.1530 0.3370 ;
        RECT 3.1510 0.3300 3.8410 0.3800 ;
        RECT 0.8870 0.2460 0.9370 0.4500 ;
        RECT 0.7350 0.2460 0.7850 0.4500 ;
        RECT 2.1030 0.3370 2.1530 0.4610 ;
        RECT 1.9510 0.3370 2.0010 0.4610 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.8640 1.7020 ;
        RECT 0.2790 1.0330 0.3290 1.6420 ;
        RECT 3.9270 0.9120 3.9770 1.6420 ;
        RECT 4.2310 0.9600 4.2810 1.6420 ;
        RECT 4.5350 1.0520 4.5850 1.6420 ;
        RECT 0.8870 1.3540 0.9370 1.6420 ;
        RECT 2.1270 1.3280 2.1770 1.6420 ;
        RECT 3.8150 1.3580 3.8650 1.6420 ;
        RECT 0.7350 1.3040 0.9370 1.3540 ;
        RECT 1.9340 1.2780 2.3360 1.3280 ;
        RECT 2.9860 1.3080 3.8650 1.3580 ;
        RECT 0.7350 1.0880 0.7850 1.3040 ;
        RECT 0.8870 1.1010 0.9370 1.3040 ;
    END
  END VDD

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7230 0.0890 3.0050 0.1390 ;
        RECT 2.9230 0.1390 3.0050 0.1750 ;
        RECT 1.7230 0.1390 1.8790 0.2180 ;
    END
    ANTENNAGATEAREA 0.0441 ;
  END RSTB

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.3590 0.6800 ;
        RECT 0.2490 0.6800 0.4210 0.7300 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.5310 0.8570 3.7030 1.0340 ;
    END
    ANTENNAGATEAREA 0.0441 ;
  END SETB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.4240 0.7250 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 4.9790 1.7730 ;
    LAYER M1 ;
      RECT 3.3030 1.2080 3.6890 1.2580 ;
      RECT 1.4790 1.2780 1.8650 1.3280 ;
      RECT 4.2880 0.6040 4.5250 0.6540 ;
      RECT 3.8150 0.7540 3.8650 1.1080 ;
      RECT 3.4550 1.1080 3.8650 1.1580 ;
      RECT 4.2880 0.5460 4.3380 0.6040 ;
      RECT 4.2880 0.6540 4.3380 0.7040 ;
      RECT 3.0140 0.5030 4.3380 0.5460 ;
      RECT 3.8150 0.7040 4.3380 0.7540 ;
      RECT 3.0140 0.4960 4.3240 0.5030 ;
      RECT 3.0140 0.5460 3.0640 0.7660 ;
      RECT 3.0140 0.7660 3.1570 0.8160 ;
      RECT 3.0140 0.4880 3.0640 0.4960 ;
      RECT 2.7110 0.4380 3.0640 0.4880 ;
      RECT 2.7110 0.4880 2.7610 1.1650 ;
      RECT 1.1910 0.2990 1.2810 0.3810 ;
      RECT 1.2150 0.3810 1.2650 0.9880 ;
      RECT 1.1910 1.0380 1.2410 1.3140 ;
      RECT 0.4310 0.9880 1.2650 1.0380 ;
      RECT 0.4310 1.0380 0.4810 1.2160 ;
      RECT 0.4310 0.8290 0.4810 0.9880 ;
      RECT 0.4310 0.5790 0.5210 0.6290 ;
      RECT 0.4310 0.4550 0.4810 0.5790 ;
      RECT 0.4310 0.7800 0.5210 0.8290 ;
      RECT 0.4710 0.6290 0.5210 0.7800 ;
      RECT 3.2430 0.1520 3.2930 0.2300 ;
      RECT 2.2950 0.2300 3.2930 0.2800 ;
      RECT 2.2950 0.2800 2.3450 0.5860 ;
      RECT 1.8590 0.5860 2.3450 0.6360 ;
      RECT 2.6190 0.1890 2.7010 0.2300 ;
      RECT 1.3430 0.6860 2.2450 0.7360 ;
      RECT 1.3430 0.7360 1.3930 1.1580 ;
      RECT 1.3430 0.4840 1.3930 0.6860 ;
      RECT 1.3430 1.2080 1.3930 1.3140 ;
      RECT 1.3430 0.3550 1.3930 0.4340 ;
      RECT 1.3430 1.1580 1.7130 1.2080 ;
      RECT 1.3430 0.4340 1.5610 0.4840 ;
      RECT 1.8590 0.7860 2.5490 0.8360 ;
      RECT 2.5590 0.6060 2.6490 0.6560 ;
      RECT 2.5990 0.6560 2.6490 1.0010 ;
      RECT 2.5590 0.4960 2.6090 0.6060 ;
      RECT 1.5500 1.0010 2.6490 1.0510 ;
      RECT 2.4070 0.4460 2.6090 0.4960 ;
      RECT 2.5590 1.0510 2.6090 1.3080 ;
      RECT 2.4070 0.3710 2.4570 0.4460 ;
      RECT 2.5590 0.3710 2.6090 0.4460 ;
      RECT 2.4070 1.3080 2.6090 1.3580 ;
      RECT 2.4070 1.2160 2.4570 1.3080 ;
      RECT 2.0860 1.1660 2.4570 1.2160 ;
      RECT 3.2070 0.6040 4.2210 0.6540 ;
      RECT 3.2070 0.6540 3.2570 0.9780 ;
      RECT 2.8460 0.9780 3.2570 1.0280 ;
      RECT 2.8460 0.5880 2.8960 0.9780 ;
      RECT 2.8460 0.5380 2.9530 0.5880 ;
      RECT 3.2260 1.4080 3.7650 1.4580 ;
      RECT 1.4190 1.4780 1.9410 1.5280 ;
      RECT 1.4190 1.5280 1.4690 1.5650 ;
      RECT 1.0990 1.5260 1.3170 1.5760 ;
      RECT 1.2670 1.4280 1.3170 1.5260 ;
      RECT 1.2670 1.3780 2.0770 1.4280 ;
      RECT 2.0270 1.4280 2.0770 1.5440 ;
      RECT 0.5830 0.6180 1.0290 0.6680 ;
      RECT 0.5830 0.6680 0.6330 0.9140 ;
      RECT 0.5830 0.4220 0.6330 0.6180 ;
      RECT 1.0390 0.5180 1.1650 0.5680 ;
      RECT 1.0390 0.3940 1.0890 0.5180 ;
      RECT 1.1150 0.5680 1.1650 0.7180 ;
      RECT 1.0390 0.7180 1.1650 0.7680 ;
      RECT 1.0390 0.7680 1.0890 0.9140 ;
      RECT 3.3450 0.7090 3.7650 0.7590 ;
      RECT 3.3450 0.7590 3.3950 1.0990 ;
      RECT 2.8350 1.0990 3.3950 1.1490 ;
      RECT 2.8350 1.1490 2.8850 1.2720 ;
      RECT 2.6590 1.2720 2.8850 1.3220 ;
      RECT 2.6590 1.3220 2.7090 1.4280 ;
      RECT 2.4670 1.4280 2.7090 1.4780 ;
      RECT 0.7950 0.0960 1.4910 0.1460 ;
      RECT 2.2860 1.5280 3.6260 1.5780 ;
    LAYER PO ;
      RECT 3.7090 1.0120 3.7390 1.6060 ;
      RECT 4.3170 0.0680 4.3470 1.6060 ;
      RECT 2.6450 0.0680 2.6750 0.6510 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 1.8850 0.7580 1.9150 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 4.7730 0.0680 4.8030 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 1.2770 0.0680 1.3070 0.5420 ;
      RECT 1.2770 0.9900 1.3070 1.6060 ;
      RECT 4.4690 0.0680 4.4990 1.6060 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 3.7090 0.0680 3.7390 0.7870 ;
      RECT 1.8850 0.0680 1.9150 0.6430 ;
      RECT 2.6450 0.8820 2.6750 1.6060 ;
      RECT 4.6210 0.0680 4.6510 1.6060 ;
  END
END DFFASRX2_LVT

MACRO DFFASX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.256 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.2560 0.0300 ;
        RECT 0.5860 0.0300 0.6360 0.1960 ;
        RECT 0.2790 0.0300 0.3290 0.4190 ;
        RECT 1.9510 0.0300 2.0010 0.4610 ;
        RECT 3.7750 0.0300 3.8250 0.2200 ;
        RECT 3.4710 0.0300 3.5210 0.3430 ;
        RECT 1.7990 0.0300 1.8490 0.3710 ;
        RECT 0.5860 0.1960 0.9370 0.2460 ;
        RECT 2.8450 0.3430 3.5370 0.3930 ;
        RECT 0.8870 0.2460 0.9370 0.4500 ;
        RECT 0.7350 0.2460 0.7850 0.4500 ;
    END
  END VSS

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.0500 1.1610 4.1600 1.2210 ;
        RECT 3.9270 1.2210 4.1600 1.2710 ;
        RECT 4.1090 0.2040 4.1590 1.1610 ;
        RECT 3.9270 1.2710 3.9770 1.5460 ;
        RECT 3.9110 0.1540 4.1590 0.2040 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.2560 1.7020 ;
        RECT 0.2790 1.0330 0.3290 1.6420 ;
        RECT 3.7750 0.9470 3.8250 1.6420 ;
        RECT 0.8870 1.3540 0.9370 1.6420 ;
        RECT 1.9750 1.3210 2.0250 1.6420 ;
        RECT 3.5110 1.3580 3.5610 1.6420 ;
        RECT 0.7350 1.3040 0.9370 1.3540 ;
        RECT 1.7740 1.2710 2.1840 1.3210 ;
        RECT 2.8340 1.3080 3.5610 1.3580 ;
        RECT 0.7350 1.0880 0.7850 1.3040 ;
        RECT 0.8870 1.1010 0.9370 1.3040 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.3590 0.6800 ;
        RECT 0.2490 0.6800 0.4210 0.7300 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2270 0.8570 3.3990 1.0340 ;
    END
    ANTENNAGATEAREA 0.0441 ;
  END SETB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.4240 0.7250 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8970 1.0090 4.0070 1.1190 ;
        RECT 3.9570 0.8540 4.0070 1.0090 ;
        RECT 3.6230 0.8040 4.0070 0.8540 ;
        RECT 3.6230 0.8540 3.6730 1.5460 ;
        RECT 3.9570 0.3590 4.0070 0.8040 ;
        RECT 3.6230 0.3090 4.0070 0.3590 ;
        RECT 3.6230 0.1480 3.6730 0.3090 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 4.3710 1.7730 ;
      RECT 2.6470 0.6640 2.9720 0.6790 ;
    LAYER M1 ;
      RECT 1.1910 0.2990 1.2810 0.3810 ;
      RECT 1.2150 0.3810 1.2650 0.9880 ;
      RECT 1.1910 1.0380 1.2410 1.3140 ;
      RECT 0.4310 0.9880 1.2650 1.0380 ;
      RECT 0.4310 1.0380 0.4810 1.2160 ;
      RECT 0.4310 0.8290 0.4810 0.9880 ;
      RECT 0.4310 0.5790 0.5210 0.6290 ;
      RECT 0.4310 0.4550 0.4810 0.5790 ;
      RECT 0.4310 0.7800 0.5210 0.8290 ;
      RECT 0.4710 0.6290 0.5210 0.7800 ;
      RECT 2.1430 0.1980 2.9890 0.2480 ;
      RECT 2.9390 0.0880 2.9890 0.1980 ;
      RECT 2.4670 0.1460 2.5490 0.1980 ;
      RECT 2.1430 0.2480 2.1930 0.5380 ;
      RECT 1.7060 0.5380 2.1930 0.5880 ;
      RECT 2.1430 0.5880 2.1930 0.5900 ;
      RECT 1.6980 0.7560 2.3970 0.8060 ;
      RECT 3.8510 0.4930 3.9010 0.7040 ;
      RECT 3.8510 0.4380 3.9010 0.4430 ;
      RECT 2.5590 0.4430 3.9010 0.4930 ;
      RECT 3.5110 0.7040 3.9010 0.7540 ;
      RECT 3.5110 0.7540 3.5610 1.1080 ;
      RECT 3.1510 1.1080 3.5610 1.1580 ;
      RECT 2.5590 0.6430 2.8530 0.6930 ;
      RECT 2.5590 0.4930 2.6090 0.6430 ;
      RECT 2.5590 0.4150 2.6090 0.4430 ;
      RECT 2.5590 0.6930 2.6090 1.1650 ;
      RECT 1.3430 0.6400 2.0930 0.6900 ;
      RECT 1.3430 0.4820 1.3930 0.6400 ;
      RECT 1.3430 0.6900 1.3930 1.1560 ;
      RECT 1.3430 0.4320 1.5610 0.4820 ;
      RECT 1.3430 1.1560 1.5610 1.2060 ;
      RECT 1.3430 0.3550 1.3930 0.4320 ;
      RECT 1.3430 1.2060 1.3930 1.3140 ;
      RECT 2.9320 0.6040 3.7650 0.6540 ;
      RECT 2.9320 0.6540 2.9820 0.9750 ;
      RECT 2.9320 0.5930 2.9820 0.6040 ;
      RECT 2.6880 0.9750 2.9820 1.0250 ;
      RECT 2.6950 0.5430 2.9820 0.5930 ;
      RECT 1.5500 1.0010 2.4970 1.0510 ;
      RECT 2.4470 0.6560 2.4970 1.0010 ;
      RECT 2.4070 1.0510 2.4570 1.3080 ;
      RECT 2.4070 0.6060 2.4970 0.6560 ;
      RECT 2.2550 1.3080 2.4570 1.3580 ;
      RECT 2.4070 0.4960 2.4570 0.6060 ;
      RECT 2.2550 1.2160 2.3050 1.3080 ;
      RECT 2.2550 0.4460 2.4570 0.4960 ;
      RECT 1.9340 1.1660 2.3050 1.2160 ;
      RECT 2.2550 0.3710 2.3050 0.4460 ;
      RECT 2.4070 0.3480 2.4570 0.4460 ;
      RECT 1.4190 1.4760 1.7890 1.5260 ;
      RECT 1.4190 1.5260 1.4690 1.5630 ;
      RECT 1.0990 1.5260 1.3170 1.5760 ;
      RECT 1.2670 1.4260 1.3170 1.5260 ;
      RECT 1.2670 1.3760 1.9250 1.4260 ;
      RECT 1.8750 1.4260 1.9250 1.5840 ;
      RECT 2.9220 1.5340 3.4610 1.5840 ;
      RECT 0.5830 0.6180 1.0290 0.6680 ;
      RECT 0.5830 0.6680 0.6330 0.9140 ;
      RECT 0.5830 0.4220 0.6330 0.6180 ;
      RECT 1.0390 0.5180 1.1650 0.5680 ;
      RECT 1.0390 0.3940 1.0890 0.5180 ;
      RECT 1.1150 0.5680 1.1650 0.7180 ;
      RECT 1.0390 0.7180 1.1650 0.7680 ;
      RECT 1.0390 0.7680 1.0890 0.9140 ;
      RECT 2.1340 1.5280 2.6820 1.5780 ;
      RECT 2.6320 1.4610 2.6820 1.5280 ;
      RECT 2.6320 1.4110 3.3090 1.4610 ;
      RECT 3.0510 0.7090 3.4610 0.7590 ;
      RECT 3.0510 0.7590 3.1010 1.0990 ;
      RECT 2.6830 1.0990 3.1010 1.1490 ;
      RECT 2.6830 1.1490 2.7330 1.2720 ;
      RECT 2.6830 1.0960 2.7330 1.0990 ;
      RECT 2.5070 1.2720 2.7330 1.3220 ;
      RECT 2.5070 1.3220 2.5570 1.4280 ;
      RECT 2.3150 1.4280 2.5570 1.4780 ;
      RECT 0.7950 0.0960 1.4910 0.1460 ;
      RECT 2.9990 1.2080 3.3850 1.2580 ;
    LAYER PO ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 3.7090 0.0680 3.7390 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 1.2770 0.0680 1.3070 0.5420 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 1.2770 0.9900 1.3070 1.6060 ;
      RECT 1.7330 0.7280 1.7630 1.6040 ;
      RECT 1.8850 0.0660 1.9150 1.6040 ;
      RECT 3.4050 0.0680 3.4350 0.7870 ;
      RECT 2.7970 0.0650 2.8270 1.6030 ;
      RECT 1.5810 0.0660 1.6110 1.6040 ;
      RECT 1.4290 0.0660 1.4590 1.6040 ;
      RECT 1.7330 0.0660 1.7630 0.6160 ;
      RECT 2.4930 0.8820 2.5230 1.6060 ;
      RECT 3.4050 1.0120 3.4350 1.6060 ;
      RECT 2.4930 0.0680 2.5230 0.6220 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
  END
END DFFASX1_LVT

MACRO DFFASX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.56 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.3530 0.0970 4.4630 0.2070 ;
        RECT 4.3950 0.2070 4.4450 0.2700 ;
        RECT 4.0790 0.2700 4.4450 0.3200 ;
        RECT 4.0790 0.1480 4.1290 0.2700 ;
        RECT 4.3950 0.3200 4.4450 0.9180 ;
        RECT 4.0790 0.9180 4.4450 0.9680 ;
        RECT 4.0790 0.9680 4.1290 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.7750 0.1480 3.8250 0.3940 ;
        RECT 3.7750 0.3940 4.3210 0.4440 ;
        RECT 4.2010 0.4440 4.3210 0.5110 ;
        RECT 4.2710 0.5110 4.3210 0.8040 ;
        RECT 3.7750 0.8040 4.3210 0.8540 ;
        RECT 3.7750 0.8540 3.8250 1.5460 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.5600 0.0300 ;
        RECT 0.5860 0.0300 0.6360 0.1960 ;
        RECT 3.6230 0.0300 3.6730 0.4080 ;
        RECT 4.2310 0.0300 4.2810 0.2200 ;
        RECT 0.2790 0.0300 0.3290 0.4190 ;
        RECT 1.9510 0.0300 2.0010 0.4610 ;
        RECT 3.9280 0.0300 3.9780 0.3120 ;
        RECT 1.7990 0.0300 1.8490 0.3710 ;
        RECT 3.4710 0.0300 3.5210 0.3430 ;
        RECT 0.5860 0.1960 0.9370 0.2460 ;
        RECT 2.8450 0.3430 3.5370 0.3930 ;
        RECT 0.8870 0.2460 0.9370 0.4500 ;
        RECT 0.7350 0.2460 0.7850 0.4500 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.5600 1.7020 ;
        RECT 0.2790 1.0330 0.3290 1.6420 ;
        RECT 3.6230 0.9120 3.6730 1.6420 ;
        RECT 3.9270 0.9600 3.9770 1.6420 ;
        RECT 4.2310 1.0520 4.2810 1.6420 ;
        RECT 0.8870 1.3540 0.9370 1.6420 ;
        RECT 1.9750 1.3210 2.0250 1.6420 ;
        RECT 3.5110 1.3580 3.5610 1.6420 ;
        RECT 0.7350 1.3040 0.9370 1.3540 ;
        RECT 1.7740 1.2710 2.1840 1.3210 ;
        RECT 2.8340 1.3080 3.5610 1.3580 ;
        RECT 0.7350 1.0880 0.7850 1.3040 ;
        RECT 0.8870 1.1010 0.9370 1.3040 ;
    END
  END VDD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.5530 0.3590 0.6800 ;
        RECT 0.2490 0.6800 0.4210 0.7300 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2270 0.8570 3.3990 1.0340 ;
    END
    ANTENNAGATEAREA 0.0441 ;
  END SETB

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.4240 0.7250 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 4.6750 1.7730 ;
      RECT 2.6600 0.6710 2.9640 0.6790 ;
    LAYER M1 ;
      RECT 1.1910 0.2990 1.2810 0.3810 ;
      RECT 1.2150 0.3810 1.2650 0.9880 ;
      RECT 1.1910 1.0380 1.2410 1.3140 ;
      RECT 0.4310 0.9880 1.2650 1.0380 ;
      RECT 0.4310 1.0380 0.4810 1.2160 ;
      RECT 0.4310 0.8290 0.4810 0.9880 ;
      RECT 0.4310 0.5790 0.5210 0.6290 ;
      RECT 0.4310 0.4550 0.4810 0.5790 ;
      RECT 0.4310 0.7800 0.5210 0.8290 ;
      RECT 0.4710 0.6290 0.5210 0.7800 ;
      RECT 2.1430 0.2300 2.9890 0.2800 ;
      RECT 2.9390 0.0880 2.9890 0.2300 ;
      RECT 2.4670 0.1780 2.5490 0.2300 ;
      RECT 2.1430 0.2800 2.1930 0.5380 ;
      RECT 1.7060 0.5380 2.1930 0.5880 ;
      RECT 2.1430 0.5880 2.1930 0.5900 ;
      RECT 1.6980 0.7560 2.3970 0.8060 ;
      RECT 3.9840 0.6040 4.2210 0.6540 ;
      RECT 3.5110 0.7540 3.5610 1.1080 ;
      RECT 3.2080 0.4930 3.2580 0.5030 ;
      RECT 3.1510 1.1080 3.5610 1.1580 ;
      RECT 2.5590 0.4430 3.2580 0.4930 ;
      RECT 3.9840 0.6540 4.0340 0.7040 ;
      RECT 3.9840 0.5530 4.0340 0.6040 ;
      RECT 3.2080 0.5030 4.0340 0.5530 ;
      RECT 3.5110 0.7040 4.0340 0.7540 ;
      RECT 2.5590 0.4930 2.6090 0.6430 ;
      RECT 2.5590 0.6430 2.8530 0.6930 ;
      RECT 2.5590 0.6930 2.6090 1.1650 ;
      RECT 1.3430 0.6400 2.0930 0.6900 ;
      RECT 1.3430 0.6900 1.3930 1.1560 ;
      RECT 1.3430 0.4820 1.3930 0.6400 ;
      RECT 1.3430 1.1560 1.5610 1.2060 ;
      RECT 1.3430 0.4320 1.5610 0.4820 ;
      RECT 1.3430 1.2060 1.3930 1.3140 ;
      RECT 1.3430 0.3550 1.3930 0.4320 ;
      RECT 2.9320 0.6040 3.9170 0.6540 ;
      RECT 2.9320 0.6540 2.9820 0.9750 ;
      RECT 2.9320 0.5930 2.9820 0.6040 ;
      RECT 2.6880 0.9750 2.9820 1.0250 ;
      RECT 2.6950 0.5440 2.9820 0.5930 ;
      RECT 2.6950 0.5430 2.9510 0.5440 ;
      RECT 2.4070 0.6060 2.4970 0.6560 ;
      RECT 2.4470 0.6560 2.4970 1.0010 ;
      RECT 2.4070 0.4960 2.4570 0.6060 ;
      RECT 1.5500 1.0010 2.4970 1.0510 ;
      RECT 2.2550 0.4460 2.4570 0.4960 ;
      RECT 2.4070 1.0510 2.4570 1.3080 ;
      RECT 2.2550 0.3710 2.3050 0.4460 ;
      RECT 2.4070 0.3710 2.4570 0.4460 ;
      RECT 2.2550 1.3080 2.4570 1.3580 ;
      RECT 2.2550 1.2160 2.3050 1.3080 ;
      RECT 1.9340 1.1660 2.3050 1.2160 ;
      RECT 1.4190 1.4760 1.7890 1.5260 ;
      RECT 1.4190 1.5260 1.4690 1.5630 ;
      RECT 3.0510 0.7090 3.4610 0.7590 ;
      RECT 3.0510 0.7590 3.1010 1.0990 ;
      RECT 2.6830 1.0990 3.1010 1.1490 ;
      RECT 2.6830 1.1490 2.7330 1.2720 ;
      RECT 2.6830 1.0960 2.7330 1.0990 ;
      RECT 2.5070 1.2720 2.7330 1.3220 ;
      RECT 2.5070 1.3220 2.5570 1.4280 ;
      RECT 2.3150 1.4280 2.5570 1.4780 ;
      RECT 1.0990 1.5260 1.3170 1.5760 ;
      RECT 1.2670 1.4260 1.3170 1.5260 ;
      RECT 1.2670 1.3760 1.9250 1.4260 ;
      RECT 1.8750 1.4260 1.9250 1.5840 ;
      RECT 2.9220 1.5340 3.4610 1.5840 ;
      RECT 0.5830 0.6180 1.0290 0.6680 ;
      RECT 0.5830 0.6680 0.6330 0.9140 ;
      RECT 0.5830 0.4220 0.6330 0.6180 ;
      RECT 1.0390 0.5180 1.1650 0.5680 ;
      RECT 1.0390 0.3940 1.0890 0.5180 ;
      RECT 1.1150 0.5680 1.1650 0.7180 ;
      RECT 1.0390 0.7180 1.1650 0.7680 ;
      RECT 1.0390 0.7680 1.0890 0.9140 ;
      RECT 2.1340 1.5280 2.6820 1.5780 ;
      RECT 2.6320 1.4610 2.6820 1.5280 ;
      RECT 2.6320 1.4110 3.3090 1.4610 ;
      RECT 0.7950 0.0960 1.4910 0.1460 ;
      RECT 2.9990 1.2080 3.3850 1.2580 ;
    LAYER PO ;
      RECT 2.4930 0.0680 2.5230 0.6220 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 1.2770 0.0680 1.3070 0.5420 ;
      RECT 3.7090 0.0680 3.7390 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 4.4690 0.0680 4.4990 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 4.3170 0.0680 4.3470 1.6060 ;
      RECT 1.2770 0.9900 1.3070 1.6060 ;
      RECT 1.7330 0.7280 1.7630 1.6040 ;
      RECT 1.8850 0.0660 1.9150 1.6040 ;
      RECT 3.4050 0.0680 3.4350 0.7870 ;
      RECT 2.7970 0.0650 2.8270 1.6030 ;
      RECT 1.5810 0.0660 1.6110 1.6040 ;
      RECT 1.4290 0.0660 1.4590 1.6040 ;
      RECT 1.7330 0.0660 1.7630 0.6160 ;
      RECT 2.4930 0.8820 2.5230 1.6060 ;
      RECT 3.4050 1.0120 3.4350 1.6060 ;
  END
END DFFASX2_LVT

MACRO BUSKP_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.824 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 1.1590 1.5850 1.2090 ;
        RECT 0.2490 0.8150 0.2990 1.1590 ;
        RECT 0.8870 1.2090 0.9370 1.4780 ;
        RECT 1.5350 0.3090 1.5850 1.1590 ;
        RECT 0.2490 0.7080 0.3590 0.8150 ;
        RECT 0.5830 0.2590 1.5850 0.3090 ;
        RECT 0.2490 0.6580 0.4210 0.7080 ;
        RECT 0.5830 0.1370 0.6330 0.2590 ;
        RECT 0.5830 0.3090 0.6330 0.3110 ;
    END
    ANTENNADIFFAREA 0.0774 ;
    ANTENNAGATEAREA 0.0774 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.8240 1.7020 ;
        RECT 0.2790 1.2880 0.3290 1.6420 ;
        RECT 0.5830 1.3180 0.6330 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.8240 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.4810 ;
        RECT 1.4950 0.0300 1.5450 0.2090 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.9390 1.7730 ;
    LAYER M1 ;
      RECT 0.5430 0.3730 1.4850 0.4230 ;
      RECT 0.5370 0.3980 0.5870 1.0990 ;
      RECT 0.4310 0.3730 0.5870 0.4230 ;
      RECT 0.4150 1.0490 0.5570 1.0990 ;
      RECT 0.4310 0.1330 0.4810 0.4910 ;
      RECT 0.4310 0.7580 0.4810 1.0740 ;
      RECT 0.4710 0.7570 0.4810 0.7580 ;
    LAYER PO ;
      RECT 1.5810 0.0730 1.6110 1.6040 ;
      RECT 1.2770 0.0730 1.3070 1.6040 ;
      RECT 1.4290 0.0730 1.4590 1.6040 ;
      RECT 1.7330 0.0730 1.7630 1.6040 ;
      RECT 1.1250 0.0730 1.1550 1.6040 ;
      RECT 0.8210 0.0730 0.8510 1.6040 ;
      RECT 0.9730 0.0730 1.0030 1.6040 ;
      RECT 0.0610 0.0730 0.0910 1.6040 ;
      RECT 0.2130 0.0730 0.2430 1.6040 ;
      RECT 0.6690 0.0730 0.6990 1.6040 ;
      RECT 0.3650 0.0730 0.3950 1.6040 ;
      RECT 0.5170 0.0730 0.5470 1.6040 ;
  END
END BUSKP_LVT

MACRO CGLNPRX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2480 1.3130 0.3590 1.4040 ;
        RECT 0.2480 1.4040 0.4210 1.4540 ;
    END
    ANTENNAGATEAREA 0.0234 ;
  END EN

  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2890 0.8340 3.4370 0.8840 ;
        RECT 3.2890 0.8840 3.3990 0.9670 ;
        RECT 3.3870 0.5850 3.4370 0.8340 ;
        RECT 3.3190 0.9670 3.3690 1.5610 ;
        RECT 3.3190 0.5350 3.4370 0.5850 ;
        RECT 3.3190 0.3140 3.3690 0.5350 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END GCLK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.8000 1.7020 ;
        RECT 3.1670 0.9260 3.2170 1.6420 ;
        RECT 1.3840 1.4760 1.4340 1.6420 ;
        RECT 3.4710 0.9260 3.5210 1.6420 ;
        RECT 2.9480 1.2540 2.9980 1.6420 ;
        RECT 0.5820 1.4260 1.4340 1.4760 ;
        RECT 1.7920 1.2040 2.9980 1.2540 ;
        RECT 0.5820 0.8260 0.6320 1.4260 ;
        RECT 1.0390 1.1520 1.0890 1.4260 ;
        RECT 0.8870 1.1650 0.9370 1.4260 ;
        RECT 2.1030 0.7580 2.1530 1.2040 ;
        RECT 2.4070 0.7580 2.4570 1.2040 ;
        RECT 1.7920 1.1020 1.8420 1.2040 ;
        RECT 2.7110 0.7560 2.7610 1.2040 ;
        RECT 1.6470 1.0520 1.8420 1.1020 ;
        RECT 1.6470 0.9280 1.6970 1.0520 ;
    END
  END VDD

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4910 0.6130 0.6630 0.6630 ;
        RECT 0.5530 0.5530 0.6630 0.6130 ;
    END
    ANTENNAGATEAREA 0.0234 ;
  END SE

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.8000 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.3370 ;
        RECT 0.5830 0.0300 0.6330 0.2820 ;
        RECT 3.5130 0.0300 3.5630 0.1970 ;
        RECT 3.0150 0.0300 3.0650 0.3210 ;
        RECT 2.7110 0.0300 2.7610 0.1900 ;
        RECT 0.5830 0.2820 1.0890 0.3320 ;
        RECT 3.4710 0.1970 3.5630 0.2470 ;
        RECT 3.0150 0.3210 3.2170 0.3710 ;
        RECT 1.6470 0.1900 2.7610 0.2400 ;
        RECT 0.8870 0.3320 0.9370 0.5320 ;
        RECT 1.0390 0.3320 1.0890 0.5460 ;
        RECT 1.0390 0.1880 1.0890 0.2820 ;
        RECT 3.4710 0.2470 3.5210 0.3710 ;
        RECT 3.1670 0.1970 3.2170 0.3210 ;
        RECT 2.4080 0.2400 2.4580 0.4400 ;
        RECT 2.1030 0.2400 2.1530 0.5320 ;
        RECT 1.6470 0.2400 1.6970 0.4080 ;
        RECT 1.6470 0.1890 1.6970 0.1900 ;
        RECT 2.7110 0.2400 2.7610 0.3480 ;
    END
  END VSS

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 0.0960 0.8770 0.2250 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 3.9150 1.7870 ;
    LAYER M1 ;
      RECT 2.5990 0.6140 3.0050 0.6640 ;
      RECT 2.5990 0.6640 2.6490 0.7550 ;
      RECT 2.5990 0.5850 2.6490 0.6140 ;
      RECT 2.5590 0.7550 2.6490 0.8050 ;
      RECT 2.5590 0.5180 2.6490 0.5850 ;
      RECT 2.5590 0.8050 2.6090 1.1130 ;
      RECT 2.5590 0.3190 2.6090 0.5180 ;
      RECT 2.2950 0.6350 2.5490 0.6850 ;
      RECT 2.2950 0.6850 2.3450 0.7550 ;
      RECT 2.2950 0.5940 2.3450 0.6350 ;
      RECT 2.2550 0.7550 2.3450 0.8050 ;
      RECT 2.2550 0.5280 2.3450 0.5940 ;
      RECT 2.2550 0.8050 2.3050 1.1130 ;
      RECT 2.2550 0.3280 2.3050 0.5280 ;
      RECT 1.6890 1.5340 2.8530 1.5840 ;
      RECT 1.1910 0.8500 1.2410 1.2100 ;
      RECT 1.1470 0.8000 1.2410 0.8500 ;
      RECT 1.1470 0.5680 1.1970 0.8000 ;
      RECT 1.1470 0.5180 1.2410 0.5680 ;
      RECT 1.1910 0.2460 1.2410 0.5180 ;
      RECT 1.1910 0.1960 1.4850 0.2460 ;
      RECT 1.6890 1.2600 1.7390 1.5340 ;
      RECT 1.1910 1.2100 1.7390 1.2600 ;
      RECT 3.2270 0.0970 3.4620 0.1470 ;
      RECT 3.1050 0.6500 3.3090 0.7000 ;
      RECT 3.1050 0.5380 3.1550 0.6500 ;
      RECT 3.1050 0.7000 3.1550 0.7140 ;
      RECT 2.8630 0.4880 3.1550 0.5380 ;
      RECT 3.0150 0.7140 3.1550 0.7640 ;
      RECT 2.8630 0.1760 2.9130 0.4880 ;
      RECT 3.0150 0.7640 3.0650 1.1170 ;
      RECT 0.9470 0.0880 1.6370 0.1380 ;
      RECT 1.9910 0.6550 2.2450 0.7050 ;
      RECT 1.4550 0.5080 1.5050 0.8860 ;
      RECT 1.4550 0.8860 1.5450 0.9360 ;
      RECT 1.4950 0.3510 1.5450 0.4580 ;
      RECT 1.4950 0.9360 1.5450 1.1200 ;
      RECT 1.9920 0.5080 2.0420 0.6550 ;
      RECT 1.9920 0.7050 2.0420 0.7690 ;
      RECT 1.4550 0.4730 2.0420 0.5080 ;
      RECT 1.9510 0.7690 2.0420 0.9330 ;
      RECT 1.9510 0.9330 2.0010 1.1020 ;
      RECT 1.9510 0.3510 2.0010 0.4580 ;
      RECT 1.4560 0.4580 2.0420 0.4730 ;
      RECT 0.7350 0.6180 1.0290 0.6680 ;
      RECT 0.7350 0.6680 0.7850 1.1900 ;
      RECT 0.7350 0.4180 0.7850 0.6180 ;
      RECT 0.4710 1.5260 1.3330 1.5760 ;
      RECT 0.2790 1.1870 0.5210 1.2370 ;
      RECT 0.4710 1.2370 0.5210 1.5260 ;
      RECT 0.2790 0.5030 0.3290 1.1870 ;
      RECT 0.2790 0.4530 0.4810 0.5030 ;
      RECT 0.4310 0.1730 0.4810 0.4530 ;
      RECT 1.5550 0.6540 1.7710 0.7040 ;
      RECT 1.7210 0.6170 1.7710 0.6540 ;
      RECT 1.7210 0.5670 1.9420 0.6170 ;
      RECT 1.2470 0.6450 1.3930 0.6950 ;
      RECT 1.3430 0.6950 1.3930 1.1600 ;
      RECT 1.3430 0.3260 1.3930 0.6450 ;
      RECT 1.4000 1.3250 1.6370 1.3750 ;
      RECT 1.7070 0.0890 2.5490 0.1390 ;
    LAYER PO ;
      RECT 3.7090 0.1080 3.7390 1.5900 ;
      RECT 2.7970 0.1080 2.8270 1.5990 ;
      RECT 3.5570 0.1080 3.5870 1.5900 ;
      RECT 3.2530 0.0860 3.2830 1.6100 ;
      RECT 1.8850 0.0690 1.9150 0.6720 ;
      RECT 1.4290 0.0670 1.4590 0.6420 ;
      RECT 1.7330 0.0720 1.7630 1.5900 ;
      RECT 1.8850 0.7720 1.9150 1.5940 ;
      RECT 3.4050 0.0860 3.4350 1.6100 ;
      RECT 2.4930 0.0730 2.5230 1.5950 ;
      RECT 2.6450 0.0740 2.6750 1.5950 ;
      RECT 3.1010 0.1090 3.1310 1.6080 ;
      RECT 0.0610 0.1090 0.0910 1.5760 ;
      RECT 0.3650 0.1070 0.3950 1.5760 ;
      RECT 0.2130 0.1090 0.2430 1.5760 ;
      RECT 1.5810 0.0650 1.6110 1.5870 ;
      RECT 1.4290 0.7420 1.4590 1.5870 ;
      RECT 0.6690 0.1070 0.6990 1.5810 ;
      RECT 1.2770 0.0680 1.3070 1.5880 ;
      RECT 0.8210 0.0840 0.8510 1.5810 ;
      RECT 0.9730 0.0680 1.0030 1.5810 ;
      RECT 1.1250 0.0680 1.1550 1.5850 ;
      RECT 2.3410 0.0720 2.3710 1.5960 ;
      RECT 0.5170 0.1070 0.5470 1.5810 ;
      RECT 2.0370 0.0690 2.0670 1.5940 ;
      RECT 2.9490 0.1080 2.9790 1.6060 ;
      RECT 2.1890 0.0700 2.2190 1.5960 ;
  END
END CGLNPRX2_LVT

MACRO CGLNPRX8_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.712 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 0.0960 0.8770 0.2250 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.7120 0.0300 ;
        RECT 3.0150 0.0300 3.0650 0.1970 ;
        RECT 0.2790 0.0300 0.3290 0.2400 ;
        RECT 0.5830 0.0300 0.6330 0.2820 ;
        RECT 2.7110 0.0300 2.7610 0.1900 ;
        RECT 3.0150 0.1970 4.4330 0.2470 ;
        RECT 0.5830 0.2820 1.0890 0.3320 ;
        RECT 1.6470 0.1900 2.7610 0.2400 ;
        RECT 4.3830 0.2470 4.4330 0.5610 ;
        RECT 3.7750 0.2470 3.8250 0.5610 ;
        RECT 4.0790 0.2470 4.1290 0.5610 ;
        RECT 3.4710 0.2470 3.5210 0.3710 ;
        RECT 3.1670 0.2470 3.2170 0.3710 ;
        RECT 3.0150 0.2470 3.0650 0.3710 ;
        RECT 1.0390 0.3320 1.0890 0.5460 ;
        RECT 1.0390 0.1880 1.0890 0.2820 ;
        RECT 0.8870 0.3320 0.9370 0.5320 ;
        RECT 2.4080 0.2400 2.4580 0.4400 ;
        RECT 2.1030 0.2400 2.1530 0.5320 ;
        RECT 1.6470 0.2400 1.6970 0.4080 ;
        RECT 1.6470 0.1890 1.6970 0.1900 ;
        RECT 2.7110 0.2400 2.7610 0.3480 ;
    END
  END VSS

  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.2890 0.8340 3.4370 0.8840 ;
        RECT 3.2890 0.8840 3.3990 0.9670 ;
        RECT 3.3870 0.7030 3.4370 0.8340 ;
        RECT 3.3190 0.9670 3.3690 1.5610 ;
        RECT 3.3870 0.6530 4.2810 0.7030 ;
        RECT 3.3870 0.5920 3.4370 0.6530 ;
        RECT 4.2310 0.7030 4.2810 1.5700 ;
        RECT 4.2310 0.3480 4.2810 0.6530 ;
        RECT 3.9270 0.7030 3.9770 1.5600 ;
        RECT 3.9270 0.3480 3.9770 0.6530 ;
        RECT 3.6230 0.7030 3.6730 1.5600 ;
        RECT 3.6230 0.3480 3.6730 0.6530 ;
        RECT 3.3190 0.5420 3.4370 0.5920 ;
        RECT 3.3190 0.3260 3.3690 0.5420 ;
    END
    ANTENNADIFFAREA 0.5952 ;
  END GCLK

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4910 0.6130 0.6630 0.6630 ;
        RECT 0.5530 0.5530 0.6630 0.6130 ;
    END
    ANTENNAGATEAREA 0.0285 ;
  END SE

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.7120 1.7020 ;
        RECT 3.7750 0.8340 3.8250 1.6420 ;
        RECT 3.1670 0.9260 3.2170 1.6420 ;
        RECT 3.4710 0.9260 3.5210 1.6420 ;
        RECT 1.3840 1.4760 1.4340 1.6420 ;
        RECT 4.0790 0.8340 4.1290 1.6420 ;
        RECT 4.3830 0.8340 4.4330 1.6420 ;
        RECT 2.9480 1.2540 2.9980 1.6420 ;
        RECT 0.5820 1.4260 1.4340 1.4760 ;
        RECT 1.7920 1.2040 2.9980 1.2540 ;
        RECT 0.5820 0.8260 0.6320 1.4260 ;
        RECT 0.8870 1.1650 0.9370 1.4260 ;
        RECT 1.0390 1.1520 1.0890 1.4260 ;
        RECT 2.1030 0.7580 2.1530 1.2040 ;
        RECT 1.7920 1.1020 1.8420 1.2040 ;
        RECT 2.4070 0.7580 2.4570 1.2040 ;
        RECT 2.7110 0.7560 2.7610 1.2040 ;
        RECT 1.6470 1.0520 1.8420 1.1020 ;
        RECT 1.6470 0.9280 1.6970 1.0520 ;
    END
  END VDD

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2480 0.4010 0.3590 0.4050 ;
        RECT 0.2480 0.4050 0.4210 0.4550 ;
        RECT 0.2480 0.4550 0.3590 0.5110 ;
    END
    ANTENNAGATEAREA 0.0285 ;
  END EN
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 4.8270 1.7860 ;
    LAYER M1 ;
      RECT 2.2950 0.6350 2.5490 0.6850 ;
      RECT 2.2950 0.6850 2.3450 0.7550 ;
      RECT 2.2950 0.5940 2.3450 0.6350 ;
      RECT 2.2550 0.7550 2.3450 0.8050 ;
      RECT 2.2550 0.5280 2.3450 0.5940 ;
      RECT 2.2550 0.8050 2.3050 1.1130 ;
      RECT 2.2550 0.3280 2.3050 0.5280 ;
      RECT 2.5990 0.6140 3.0050 0.6640 ;
      RECT 2.5990 0.6640 2.6490 0.7550 ;
      RECT 2.5990 0.5850 2.6490 0.6140 ;
      RECT 2.5590 0.7550 2.6490 0.8050 ;
      RECT 2.5590 0.5180 2.6490 0.5850 ;
      RECT 2.5590 0.8050 2.6090 1.1130 ;
      RECT 2.5590 0.3190 2.6090 0.5180 ;
      RECT 1.9910 0.6550 2.2450 0.7050 ;
      RECT 1.4550 0.5080 1.5050 0.8860 ;
      RECT 1.4550 0.8860 1.5450 0.9360 ;
      RECT 1.4950 0.3510 1.5450 0.4580 ;
      RECT 1.4950 0.9360 1.5450 1.1200 ;
      RECT 1.9920 0.5080 2.0420 0.6550 ;
      RECT 1.9920 0.7050 2.0420 0.7690 ;
      RECT 1.4550 0.4730 2.0420 0.5080 ;
      RECT 1.9510 0.7690 2.0420 0.9330 ;
      RECT 1.9510 0.9330 2.0010 1.1020 ;
      RECT 1.9510 0.3510 2.0010 0.4580 ;
      RECT 1.4560 0.4580 2.0420 0.4730 ;
      RECT 1.6890 1.5340 2.8530 1.5840 ;
      RECT 1.1910 0.8500 1.2410 1.2100 ;
      RECT 1.1470 0.8000 1.2410 0.8500 ;
      RECT 1.1470 0.5680 1.1970 0.8000 ;
      RECT 1.1470 0.5180 1.2410 0.5680 ;
      RECT 1.1910 0.2460 1.2410 0.5180 ;
      RECT 1.1910 0.1960 1.4850 0.2460 ;
      RECT 1.6890 1.2600 1.7390 1.5340 ;
      RECT 1.1910 1.2100 1.7390 1.2600 ;
      RECT 3.1050 0.6570 3.3090 0.7070 ;
      RECT 3.1050 0.5380 3.1550 0.6570 ;
      RECT 3.1050 0.7070 3.1550 0.7140 ;
      RECT 2.8630 0.4880 3.1550 0.5380 ;
      RECT 3.0150 0.7140 3.1550 0.7640 ;
      RECT 2.8630 0.1800 2.9130 0.4880 ;
      RECT 3.0150 0.7640 3.0650 1.1170 ;
      RECT 0.4710 1.5260 1.3330 1.5760 ;
      RECT 0.4710 1.2370 0.5210 1.5260 ;
      RECT 0.2790 1.1870 0.5210 1.2370 ;
      RECT 0.2790 0.7760 0.3290 1.1870 ;
      RECT 0.1480 0.7260 0.3290 0.7760 ;
      RECT 0.4310 0.1630 0.4810 0.2900 ;
      RECT 0.1480 0.2900 0.4810 0.3400 ;
      RECT 0.1480 0.3400 0.1980 0.7260 ;
      RECT 0.7350 0.6180 1.0290 0.6680 ;
      RECT 0.7350 0.6680 0.7850 1.1900 ;
      RECT 0.7350 0.4180 0.7850 0.6180 ;
      RECT 0.9470 0.0880 1.6370 0.1380 ;
      RECT 3.2270 0.0970 4.3730 0.1470 ;
      RECT 1.7070 0.0890 2.5490 0.1390 ;
      RECT 1.3430 0.6950 1.3930 1.1600 ;
      RECT 1.2470 0.6450 1.3930 0.6950 ;
      RECT 1.3430 0.3260 1.3930 0.6450 ;
      RECT 1.4000 1.3250 1.6370 1.3750 ;
      RECT 1.5550 0.6540 1.7710 0.7040 ;
      RECT 1.7210 0.6170 1.7710 0.6540 ;
      RECT 1.7210 0.5670 1.9420 0.6170 ;
    LAYER PO ;
      RECT 3.5570 0.0860 3.5870 1.6100 ;
      RECT 3.2530 0.0860 3.2830 1.6100 ;
      RECT 4.1650 0.0860 4.1950 1.6100 ;
      RECT 1.8850 0.7720 1.9150 1.6150 ;
      RECT 1.7330 0.0710 1.7630 1.5900 ;
      RECT 1.4290 0.0670 1.4590 0.6420 ;
      RECT 1.8850 0.0670 1.9150 0.6720 ;
      RECT 3.4050 0.0860 3.4350 1.6100 ;
      RECT 2.7970 0.1070 2.8270 1.5960 ;
      RECT 3.8610 0.0860 3.8910 1.6100 ;
      RECT 4.3170 0.0860 4.3470 1.6100 ;
      RECT 2.1890 0.0750 2.2190 1.5990 ;
      RECT 2.9490 0.1070 2.9790 1.6060 ;
      RECT 3.7090 0.0860 3.7390 1.6100 ;
      RECT 2.0370 0.0750 2.0670 1.5990 ;
      RECT 4.0130 0.0860 4.0430 1.6100 ;
      RECT 0.5170 0.1080 0.5470 1.6060 ;
      RECT 2.3410 0.0520 2.3710 1.5990 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 0.8210 0.0830 0.8510 1.6060 ;
      RECT 1.2770 0.0680 1.3070 1.6060 ;
      RECT 0.6690 0.1080 0.6990 1.6060 ;
      RECT 1.4290 0.7420 1.4590 1.5900 ;
      RECT 1.5810 0.0670 1.6110 1.5900 ;
      RECT 0.2130 0.1100 0.2430 1.6060 ;
      RECT 0.3650 0.1080 0.3950 1.6060 ;
      RECT 0.0610 0.1100 0.0910 1.6060 ;
      RECT 3.1010 0.1060 3.1310 1.6080 ;
      RECT 2.6450 0.0710 2.6750 1.5990 ;
      RECT 2.4930 0.0690 2.5230 1.5990 ;
      RECT 4.6210 0.0840 4.6510 1.5900 ;
      RECT 4.4690 0.0840 4.4990 1.5900 ;
  END
END CGLNPRX8_LVT

MACRO CGLNPSX16_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.144 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 0.8570 0.9670 0.9670 ;
        RECT 0.9170 0.6680 0.9670 0.8570 ;
        RECT 0.9170 0.6180 1.0290 0.6680 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END EN

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.3310 0.6480 2.3810 1.0090 ;
        RECT 2.2250 1.0090 2.3810 1.1190 ;
    END
    ANTENNAGATEAREA 0.027 ;
  END SE

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 7.1440 1.7020 ;
        RECT 4.8390 0.9040 4.8890 1.6420 ;
        RECT 5.1430 0.9040 5.1930 1.6420 ;
        RECT 5.4470 0.9040 5.4970 1.6420 ;
        RECT 4.5350 0.9040 4.5850 1.6420 ;
        RECT 3.7750 0.9040 3.8250 1.6420 ;
        RECT 4.0790 0.9040 4.1290 1.6420 ;
        RECT 3.3190 0.9040 3.3690 1.6420 ;
        RECT 6.0550 0.9040 6.1050 1.6420 ;
        RECT 6.3590 0.9040 6.4090 1.6420 ;
        RECT 6.6630 0.9040 6.7130 1.6420 ;
        RECT 5.7510 0.9040 5.8010 1.6420 ;
        RECT 0.5430 1.3540 0.5930 1.6420 ;
        RECT 2.7110 1.3660 2.7610 1.6420 ;
        RECT 0.4310 1.3040 1.5450 1.3540 ;
        RECT 2.0870 1.3160 2.7610 1.3660 ;
        RECT 0.4310 1.0880 0.4810 1.3040 ;
        RECT 0.5830 0.9490 0.6330 1.3040 ;
        RECT 1.4950 0.7500 1.5450 1.3040 ;
        RECT 0.8870 1.0370 0.9370 1.3040 ;
        RECT 2.7110 1.0920 2.7610 1.3160 ;
    END
  END VDD

  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.7850 1.1610 6.9050 1.2710 ;
        RECT 6.8150 1.2710 6.8650 1.5460 ;
        RECT 6.8550 0.8540 6.9050 1.1610 ;
        RECT 4.3830 0.8040 6.9050 0.8540 ;
        RECT 6.5110 0.8540 6.5610 1.5460 ;
        RECT 6.2070 0.8540 6.2570 1.5460 ;
        RECT 5.9030 0.8540 5.9530 1.5460 ;
        RECT 5.5990 0.8540 5.6490 1.5460 ;
        RECT 5.2950 0.8540 5.3450 1.5460 ;
        RECT 4.9910 0.8540 5.0410 1.5460 ;
        RECT 4.6870 0.8540 4.7370 1.5460 ;
        RECT 4.3830 0.8540 4.4330 1.5460 ;
        RECT 6.8550 0.5540 6.9050 0.8040 ;
        RECT 4.3830 0.5040 6.9050 0.5540 ;
        RECT 6.8150 0.1480 6.8650 0.5040 ;
        RECT 6.5110 0.1480 6.5610 0.5040 ;
        RECT 6.2070 0.1480 6.2570 0.5040 ;
        RECT 5.9030 0.1480 5.9530 0.5040 ;
        RECT 5.5990 0.1480 5.6490 0.5040 ;
        RECT 5.2950 0.1480 5.3450 0.5040 ;
        RECT 4.9910 0.1480 5.0410 0.5040 ;
        RECT 4.6870 0.1480 4.7370 0.5040 ;
        RECT 4.3830 0.1480 4.4330 0.5040 ;
    END
    ANTENNADIFFAREA 1.2904 ;
  END GCLK

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 7.1440 0.0300 ;
        RECT 4.8390 0.0300 4.8890 0.4540 ;
        RECT 5.1430 0.0300 5.1930 0.4540 ;
        RECT 5.4470 0.0300 5.4970 0.4540 ;
        RECT 4.5350 0.0300 4.5850 0.4540 ;
        RECT 3.7750 0.0300 3.8250 0.4540 ;
        RECT 4.0790 0.0300 4.1290 0.4540 ;
        RECT 3.3190 0.0300 3.3690 0.4540 ;
        RECT 5.7510 0.0300 5.8010 0.4540 ;
        RECT 6.0550 0.0300 6.1050 0.4540 ;
        RECT 6.3590 0.0300 6.4090 0.4540 ;
        RECT 6.6630 0.0300 6.7130 0.4540 ;
        RECT 0.4310 0.0300 0.4810 0.1960 ;
        RECT 2.9030 0.0300 2.9530 0.1960 ;
        RECT 0.4310 0.1960 0.9370 0.2460 ;
        RECT 2.4070 0.1960 2.9530 0.2460 ;
        RECT 0.4310 0.2460 0.4810 0.4500 ;
        RECT 0.8870 0.2460 0.9370 0.4500 ;
        RECT 0.5830 0.2460 0.6330 0.4500 ;
        RECT 2.8630 0.2460 2.9130 0.4670 ;
        RECT 2.4070 0.2460 2.4570 0.3180 ;
        RECT 1.4790 0.3180 2.4570 0.3680 ;
        RECT 2.4070 0.3680 2.4570 0.4720 ;
    END
  END VSS

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 1.4240 0.4210 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 7.2590 1.7870 ;
    LAYER M1 ;
      RECT 4.2710 0.6040 6.8050 0.6540 ;
      RECT 3.6230 0.1480 3.6730 0.5040 ;
      RECT 3.6230 0.8540 3.6730 1.5460 ;
      RECT 3.9270 0.1480 3.9770 0.5040 ;
      RECT 3.9270 0.8540 3.9770 1.5460 ;
      RECT 4.2310 0.1480 4.2810 0.5040 ;
      RECT 4.2710 0.5540 4.3210 0.6040 ;
      RECT 4.2710 0.6540 4.3210 0.8040 ;
      RECT 4.2310 0.8540 4.2810 1.5460 ;
      RECT 3.6230 0.8040 4.3210 0.8540 ;
      RECT 3.6230 0.5040 4.3210 0.5540 ;
      RECT 3.5110 0.6040 4.2210 0.6540 ;
      RECT 3.1670 0.8540 3.2170 1.5460 ;
      RECT 3.1670 0.1480 3.2170 0.5040 ;
      RECT 3.5110 0.6540 3.5610 0.8040 ;
      RECT 3.5110 0.5540 3.5610 0.6040 ;
      RECT 3.4710 0.8540 3.5210 1.5460 ;
      RECT 3.4710 0.1480 3.5210 0.5040 ;
      RECT 3.1670 0.8040 3.5610 0.8540 ;
      RECT 3.1670 0.5040 3.5610 0.5540 ;
      RECT 2.5590 0.6300 3.0050 0.6800 ;
      RECT 2.2550 0.5720 2.3050 0.5920 ;
      RECT 2.2550 0.5020 2.3050 0.5220 ;
      RECT 2.5590 0.6800 2.6090 1.2660 ;
      RECT 2.5590 0.5720 2.6090 0.6300 ;
      RECT 2.5590 0.4790 2.6090 0.5220 ;
      RECT 2.2550 0.5220 2.6090 0.5720 ;
      RECT 3.0550 0.6040 3.4610 0.6540 ;
      RECT 3.0550 0.6540 3.1050 0.8860 ;
      RECT 3.0550 0.5670 3.1050 0.6040 ;
      RECT 3.0150 0.8860 3.1050 0.9360 ;
      RECT 2.6940 0.5170 3.1050 0.5670 ;
      RECT 3.0150 0.9360 3.0650 1.3580 ;
      RECT 0.2790 0.6180 0.7250 0.6680 ;
      RECT 0.2790 0.6680 0.3290 0.9140 ;
      RECT 0.2790 0.4220 0.3290 0.6180 ;
      RECT 0.7350 0.5180 0.8610 0.5680 ;
      RECT 0.8110 0.5680 0.8610 0.7180 ;
      RECT 0.7350 0.7180 0.8610 0.7680 ;
      RECT 0.7350 0.3940 0.7850 0.5180 ;
      RECT 0.7350 0.7680 0.7850 0.9140 ;
      RECT 1.6470 0.7510 1.7370 0.8010 ;
      RECT 1.6470 0.8010 1.6970 0.9920 ;
      RECT 1.6870 0.6680 1.7370 0.7510 ;
      RECT 1.6870 0.6180 2.0930 0.6680 ;
      RECT 1.6870 0.5680 1.7370 0.6180 ;
      RECT 1.6310 0.5180 1.7370 0.5680 ;
      RECT 1.6070 1.0420 1.9250 1.0920 ;
      RECT 1.8750 0.7180 1.9250 1.0420 ;
      RECT 1.6070 1.0920 1.6570 1.5260 ;
      RECT 0.6430 1.5260 1.6570 1.5760 ;
      RECT 1.7070 1.5310 1.9450 1.5810 ;
      RECT 1.9750 0.7280 2.1930 0.7780 ;
      RECT 2.1430 0.4680 2.1930 0.7280 ;
      RECT 1.9750 0.7780 2.0250 1.2200 ;
      RECT 1.7830 1.2200 2.0250 1.2700 ;
      RECT 1.3430 0.6180 1.6370 0.6680 ;
      RECT 1.3430 0.4180 2.1930 0.4680 ;
      RECT 1.3430 0.2820 1.3930 0.4180 ;
      RECT 1.3430 0.4680 1.3930 0.6180 ;
      RECT 1.3430 0.6680 1.3930 1.2540 ;
      RECT 1.0390 1.2040 1.2410 1.2540 ;
      RECT 1.0390 0.7500 1.0890 1.2040 ;
      RECT 1.1910 0.5680 1.2410 1.2040 ;
      RECT 1.0390 0.1960 1.0890 0.5180 ;
      RECT 1.1910 0.2820 1.2410 0.5180 ;
      RECT 1.0390 0.5180 1.2410 0.5680 ;
      RECT 2.0110 1.5310 2.5490 1.5810 ;
      RECT 0.6430 0.0960 2.8530 0.1460 ;
    LAYER PO ;
      RECT 1.8850 0.0680 1.9150 0.8120 ;
      RECT 4.7730 0.0680 4.8030 1.6060 ;
      RECT 5.3810 0.0680 5.4110 1.6060 ;
      RECT 5.8370 0.0680 5.8670 1.6060 ;
      RECT 5.5330 0.0680 5.5630 1.6060 ;
      RECT 4.9250 0.0680 4.9550 1.6060 ;
      RECT 5.2290 0.0680 5.2590 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 5.0770 0.0680 5.1070 1.6060 ;
      RECT 5.6850 0.0680 5.7150 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 3.7090 0.0680 3.7390 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 4.3170 0.0680 4.3470 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 6.2930 0.0680 6.3230 1.6060 ;
      RECT 5.9890 0.0680 6.0190 1.6060 ;
      RECT 6.1410 0.0680 6.1710 1.6060 ;
      RECT 6.4450 0.0680 6.4750 1.6060 ;
      RECT 6.5970 0.0680 6.6270 1.6060 ;
      RECT 7.0530 0.0680 7.0830 1.6060 ;
      RECT 6.7490 0.0680 6.7790 1.6060 ;
      RECT 6.9010 0.0680 6.9310 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 1.8850 1.0820 1.9150 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 4.6210 0.0680 4.6510 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 4.4690 0.0680 4.4990 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 1.2770 0.0680 1.3070 0.6420 ;
      RECT 1.2770 0.9900 1.3070 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
  END
END CGLNPSX16_LVT

MACRO CGLNPSX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 0.8570 0.9670 0.9670 ;
        RECT 0.9170 0.6680 0.9670 0.8570 ;
        RECT 0.9170 0.6180 1.0290 0.6680 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END EN

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2250 1.0090 2.3350 1.1190 ;
        RECT 2.2850 0.7520 2.3350 1.0090 ;
        RECT 2.2850 0.7020 2.3970 0.7520 ;
    END
    ANTENNAGATEAREA 0.0234 ;
  END SE

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.8000 1.7020 ;
        RECT 3.3190 0.9040 3.3690 1.6420 ;
        RECT 0.5430 1.3540 0.5930 1.6420 ;
        RECT 2.7110 1.3660 2.7610 1.6420 ;
        RECT 0.4310 1.3040 1.5450 1.3540 ;
        RECT 2.0870 1.3160 2.7610 1.3660 ;
        RECT 0.4310 1.0880 0.4810 1.3040 ;
        RECT 0.5830 0.9490 0.6330 1.3040 ;
        RECT 1.4950 0.7500 1.5450 1.3040 ;
        RECT 0.8870 1.0370 0.9370 1.3040 ;
        RECT 2.7110 1.0920 2.7610 1.3160 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.8000 0.0300 ;
        RECT 3.3190 0.0300 3.3690 0.4540 ;
        RECT 0.4310 0.0300 0.4810 0.1960 ;
        RECT 2.9030 0.0300 2.9530 0.1960 ;
        RECT 0.4310 0.1960 0.9370 0.2460 ;
        RECT 2.4070 0.1960 2.9530 0.2460 ;
        RECT 0.4310 0.2460 0.4810 0.4500 ;
        RECT 0.8870 0.2460 0.9370 0.4700 ;
        RECT 0.5830 0.2460 0.6330 0.4500 ;
        RECT 2.8630 0.2460 2.9130 0.4770 ;
        RECT 2.4070 0.2460 2.4570 0.3180 ;
        RECT 1.4790 0.3180 2.4570 0.3680 ;
        RECT 2.4070 0.3680 2.4570 0.4920 ;
    END
  END VSS

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 1.4240 0.4210 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4410 1.1610 3.5610 1.2710 ;
        RECT 3.4710 1.2710 3.5210 1.5460 ;
        RECT 3.5110 0.8540 3.5610 1.1610 ;
        RECT 3.1670 0.8040 3.5610 0.8540 ;
        RECT 3.1670 0.8540 3.2170 1.5460 ;
        RECT 3.5110 0.5540 3.5610 0.8040 ;
        RECT 3.1670 0.5040 3.5610 0.5540 ;
        RECT 3.4710 0.1480 3.5210 0.5040 ;
        RECT 3.1670 0.1480 3.2170 0.5040 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END GCLK
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 3.9150 1.7870 ;
    LAYER M1 ;
      RECT 2.5590 0.6900 3.0050 0.7400 ;
      RECT 2.2550 0.4180 2.3050 0.5420 ;
      RECT 2.5590 0.7400 2.6090 1.2660 ;
      RECT 2.5590 0.5920 2.6090 0.6900 ;
      RECT 2.5590 0.3750 2.6090 0.5420 ;
      RECT 2.2550 0.5420 2.6090 0.5920 ;
      RECT 2.1430 0.4680 2.1930 0.7280 ;
      RECT 1.9750 0.7280 2.1930 0.7780 ;
      RECT 1.3430 0.6180 1.6370 0.6680 ;
      RECT 1.9750 0.7780 2.0250 1.2200 ;
      RECT 1.7830 1.2200 2.0250 1.2700 ;
      RECT 1.3430 0.4180 2.1930 0.4680 ;
      RECT 1.3430 0.4680 1.3930 0.6180 ;
      RECT 1.3430 0.2820 1.3930 0.4180 ;
      RECT 1.3430 0.6680 1.3930 1.2540 ;
      RECT 1.1910 0.2820 1.2410 0.5180 ;
      RECT 1.0390 0.1960 1.0890 0.5180 ;
      RECT 1.1910 0.5680 1.2410 1.2040 ;
      RECT 1.0390 1.2040 1.2410 1.2540 ;
      RECT 1.0390 0.7500 1.0890 1.2040 ;
      RECT 1.0390 0.5180 1.2410 0.5680 ;
      RECT 0.8110 0.5680 0.8610 0.7180 ;
      RECT 0.7350 0.7180 0.8610 0.7680 ;
      RECT 0.7350 0.5200 0.8610 0.5680 ;
      RECT 0.7350 0.5180 0.8370 0.5200 ;
      RECT 0.7350 0.3940 0.7850 0.5180 ;
      RECT 0.7350 0.7680 0.7850 0.9140 ;
      RECT 1.6070 1.0420 1.9250 1.0920 ;
      RECT 1.8750 0.7180 1.9250 1.0420 ;
      RECT 1.6070 1.0920 1.6570 1.5260 ;
      RECT 0.6430 1.5260 1.6570 1.5760 ;
      RECT 1.7070 1.5310 1.9450 1.5810 ;
      RECT 3.0550 0.6040 3.4610 0.6540 ;
      RECT 2.7110 0.4890 2.7610 0.5540 ;
      RECT 3.0550 0.6540 3.1050 0.8860 ;
      RECT 2.6940 0.5540 3.1050 0.6040 ;
      RECT 3.0150 0.8860 3.1050 0.9360 ;
      RECT 3.0150 0.5430 3.1050 0.5540 ;
      RECT 3.0150 0.9360 3.0650 1.3580 ;
      RECT 3.0150 0.2820 3.0650 0.5430 ;
      RECT 1.6470 0.7510 1.7370 0.8010 ;
      RECT 1.6470 0.8010 1.6970 0.9920 ;
      RECT 1.6870 0.6680 1.7370 0.7510 ;
      RECT 1.6870 0.6180 2.0930 0.6680 ;
      RECT 1.6870 0.5680 1.7370 0.6180 ;
      RECT 1.6310 0.5180 1.7370 0.5680 ;
      RECT 0.2790 0.6180 0.7250 0.6680 ;
      RECT 0.2790 0.6680 0.3290 0.9140 ;
      RECT 0.2790 0.4220 0.3290 0.6180 ;
      RECT 2.0110 1.5310 2.5490 1.5810 ;
      RECT 0.6430 0.0960 2.8530 0.1460 ;
    LAYER PO ;
      RECT 1.8850 0.0680 1.9150 0.8120 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 1.8850 1.0820 1.9150 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 1.2770 0.0680 1.3070 0.6420 ;
      RECT 3.7090 0.0680 3.7390 1.6060 ;
      RECT 1.2770 0.9900 1.3070 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
  END
END CGLNPSX2_LVT

MACRO CGLNPSX4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.104 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 0.8570 0.9670 0.9670 ;
        RECT 0.9170 0.6680 0.9670 0.8570 ;
        RECT 0.9170 0.6180 1.0290 0.6680 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END EN

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2250 1.0090 2.3350 1.1190 ;
        RECT 2.2850 0.7430 2.3350 1.0090 ;
        RECT 2.2850 0.6930 2.3970 0.7430 ;
    END
    ANTENNAGATEAREA 0.0234 ;
  END SE

  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.7450 1.1610 3.8650 1.2710 ;
        RECT 3.7750 1.2710 3.8250 1.5460 ;
        RECT 3.8150 0.8540 3.8650 1.1610 ;
        RECT 3.1670 0.8040 3.8650 0.8540 ;
        RECT 3.4710 0.8540 3.5210 1.5460 ;
        RECT 3.1670 0.8540 3.2170 1.5460 ;
        RECT 3.8150 0.5540 3.8650 0.8040 ;
        RECT 3.1670 0.5040 3.8650 0.5540 ;
        RECT 3.7750 0.1480 3.8250 0.5040 ;
        RECT 3.4710 0.1480 3.5210 0.5040 ;
        RECT 3.1670 0.1480 3.2170 0.5040 ;
    END
    ANTENNADIFFAREA 0.3976 ;
  END GCLK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.1040 1.7020 ;
        RECT 3.6230 0.9040 3.6730 1.6420 ;
        RECT 3.3190 0.9040 3.3690 1.6420 ;
        RECT 0.5430 1.3540 0.5930 1.6420 ;
        RECT 2.7110 1.3660 2.7610 1.6420 ;
        RECT 0.4310 1.3040 1.5450 1.3540 ;
        RECT 2.0870 1.3160 2.7610 1.3660 ;
        RECT 0.4310 1.0880 0.4810 1.3040 ;
        RECT 0.5830 0.9490 0.6330 1.3040 ;
        RECT 1.4950 0.7500 1.5450 1.3040 ;
        RECT 0.8870 1.0370 0.9370 1.3040 ;
        RECT 2.7110 1.0920 2.7610 1.3160 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.1040 0.0300 ;
        RECT 3.6230 0.0300 3.6730 0.4540 ;
        RECT 3.3190 0.0300 3.3690 0.4540 ;
        RECT 0.4310 0.0300 0.4810 0.1960 ;
        RECT 2.9030 0.0300 2.9530 0.1960 ;
        RECT 0.4310 0.1960 0.9370 0.2460 ;
        RECT 2.4070 0.1960 2.9530 0.2460 ;
        RECT 0.4310 0.2460 0.4810 0.4500 ;
        RECT 0.8870 0.2460 0.9370 0.4500 ;
        RECT 0.5830 0.2460 0.6330 0.4500 ;
        RECT 2.8630 0.2460 2.9130 0.4830 ;
        RECT 2.4070 0.2460 2.4570 0.3180 ;
        RECT 1.4790 0.3180 2.4570 0.3680 ;
        RECT 2.4070 0.3680 2.4570 0.4910 ;
    END
  END VSS

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 1.4240 0.4210 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 4.2190 1.7870 ;
    LAYER M1 ;
      RECT 2.5590 0.6920 3.0050 0.7420 ;
      RECT 2.2550 0.4180 2.3050 0.5420 ;
      RECT 2.5590 0.7420 2.6090 1.2660 ;
      RECT 2.5590 0.5920 2.6090 0.6920 ;
      RECT 2.2550 0.5420 2.6090 0.5920 ;
      RECT 2.5590 0.3810 2.6090 0.5420 ;
      RECT 0.2790 0.6180 0.7250 0.6680 ;
      RECT 0.2790 0.6680 0.3290 0.9140 ;
      RECT 0.2790 0.4220 0.3290 0.6180 ;
      RECT 0.7350 0.5180 0.8610 0.5680 ;
      RECT 0.8110 0.5680 0.8610 0.7180 ;
      RECT 0.7350 0.7180 0.8610 0.7680 ;
      RECT 0.7350 0.3940 0.7850 0.5180 ;
      RECT 0.7350 0.7680 0.7850 0.9140 ;
      RECT 1.6470 0.7510 1.7370 0.8010 ;
      RECT 1.6470 0.8010 1.6970 0.9920 ;
      RECT 1.6870 0.6680 1.7370 0.7510 ;
      RECT 1.6870 0.6180 2.0930 0.6680 ;
      RECT 1.6870 0.5680 1.7370 0.6180 ;
      RECT 1.6310 0.5180 1.7370 0.5680 ;
      RECT 3.0550 0.6210 3.7650 0.6540 ;
      RECT 2.6940 0.6040 3.7650 0.6210 ;
      RECT 2.7110 0.4970 2.7610 0.5710 ;
      RECT 3.0550 0.6540 3.1050 0.8860 ;
      RECT 2.6940 0.5710 3.1050 0.6040 ;
      RECT 3.0150 0.8860 3.1050 0.9360 ;
      RECT 3.0150 0.5540 3.1050 0.5710 ;
      RECT 3.0150 0.9360 3.0650 1.3580 ;
      RECT 3.0150 0.2820 3.0650 0.5540 ;
      RECT 2.1430 0.4680 2.1930 0.7280 ;
      RECT 1.9750 0.7280 2.1930 0.7780 ;
      RECT 1.3430 0.6180 1.6370 0.6680 ;
      RECT 1.9750 0.7780 2.0250 1.2200 ;
      RECT 1.7830 1.2200 2.0250 1.2700 ;
      RECT 1.3430 0.4180 2.1930 0.4680 ;
      RECT 1.3430 0.4680 1.3930 0.6180 ;
      RECT 1.3430 0.2820 1.3930 0.4180 ;
      RECT 1.3430 0.6680 1.3930 1.2540 ;
      RECT 1.1910 0.2820 1.2410 0.5180 ;
      RECT 1.0390 0.1960 1.0890 0.5180 ;
      RECT 1.1910 0.5680 1.2410 1.2040 ;
      RECT 1.0390 1.2040 1.2410 1.2540 ;
      RECT 1.0390 0.7500 1.0890 1.2040 ;
      RECT 1.0390 0.5180 1.2410 0.5680 ;
      RECT 1.6070 1.0420 1.9250 1.0920 ;
      RECT 1.8750 0.7180 1.9250 1.0420 ;
      RECT 1.6070 1.0920 1.6570 1.5260 ;
      RECT 0.6430 1.5260 1.6570 1.5760 ;
      RECT 1.7070 1.5310 1.9450 1.5810 ;
      RECT 2.0110 1.5310 2.5490 1.5810 ;
      RECT 0.6430 0.0960 2.8530 0.1460 ;
    LAYER PO ;
      RECT 1.8850 0.0680 1.9150 0.8120 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 1.8850 1.0820 1.9150 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 3.7090 0.0680 3.7390 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 1.2770 0.0680 1.3070 0.6420 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 1.2770 0.9900 1.3070 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
  END
END CGLNPSX4_LVT

MACRO CGLNPSX8_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.712 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 0.8570 0.9670 0.9670 ;
        RECT 0.9170 0.6680 0.9670 0.8570 ;
        RECT 0.9170 0.6180 1.0290 0.6680 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END EN

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2250 1.0090 2.3350 1.1190 ;
        RECT 2.2850 0.6990 2.3350 1.0090 ;
        RECT 2.2830 0.6490 2.3970 0.6990 ;
    END
    ANTENNAGATEAREA 0.027 ;
  END SE

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.7120 1.7020 ;
        RECT 3.3190 0.9040 3.3690 1.6420 ;
        RECT 3.6230 0.9040 3.6730 1.6420 ;
        RECT 3.9270 0.9040 3.9770 1.6420 ;
        RECT 4.2310 0.9040 4.2810 1.6420 ;
        RECT 0.5430 1.3540 0.5930 1.6420 ;
        RECT 2.7110 1.3660 2.7610 1.6420 ;
        RECT 0.4310 1.3040 1.5450 1.3540 ;
        RECT 2.0870 1.3160 2.7610 1.3660 ;
        RECT 0.4310 1.0880 0.4810 1.3040 ;
        RECT 0.5830 0.9490 0.6330 1.3040 ;
        RECT 1.4950 0.7500 1.5450 1.3040 ;
        RECT 0.8870 1.0370 0.9370 1.3040 ;
        RECT 2.7110 1.0920 2.7610 1.3160 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.7120 0.0300 ;
        RECT 3.6230 0.0300 3.6730 0.4540 ;
        RECT 3.9270 0.0300 3.9770 0.4540 ;
        RECT 4.2310 0.0300 4.2810 0.4540 ;
        RECT 3.3190 0.0300 3.3690 0.4540 ;
        RECT 0.4310 0.0300 0.4810 0.1960 ;
        RECT 2.9030 0.0300 2.9530 0.1960 ;
        RECT 0.4310 0.1960 0.9370 0.2460 ;
        RECT 2.4070 0.1960 2.9530 0.2460 ;
        RECT 0.4310 0.2460 0.4810 0.4500 ;
        RECT 0.8870 0.2460 0.9370 0.4500 ;
        RECT 0.5830 0.2460 0.6330 0.4500 ;
        RECT 2.8630 0.2460 2.9130 0.4630 ;
        RECT 2.4070 0.2460 2.4570 0.3180 ;
        RECT 1.4790 0.3180 2.4570 0.3680 ;
        RECT 2.4070 0.3680 2.4570 0.4770 ;
    END
  END VSS

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 1.4240 0.4210 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.3530 1.1610 4.4730 1.2710 ;
        RECT 4.3830 1.2710 4.4330 1.5460 ;
        RECT 4.4230 0.8540 4.4730 1.1610 ;
        RECT 3.1670 0.8040 4.4730 0.8540 ;
        RECT 4.0790 0.8540 4.1290 1.5460 ;
        RECT 3.7750 0.8540 3.8250 1.5460 ;
        RECT 3.4710 0.8540 3.5210 1.5460 ;
        RECT 3.1670 0.8540 3.2170 1.5460 ;
        RECT 4.4230 0.5540 4.4730 0.8040 ;
        RECT 3.1670 0.5040 4.4730 0.5540 ;
        RECT 4.3830 0.1480 4.4330 0.5040 ;
        RECT 4.0790 0.1480 4.1290 0.5040 ;
        RECT 3.7750 0.1480 3.8250 0.5040 ;
        RECT 3.4710 0.1480 3.5210 0.5040 ;
        RECT 3.1670 0.1480 3.2170 0.5040 ;
    END
    ANTENNADIFFAREA 0.6952 ;
  END GCLK
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 4.8270 1.7870 ;
    LAYER M1 ;
      RECT 2.5590 0.6500 3.0050 0.7000 ;
      RECT 2.2550 0.4180 2.3050 0.5420 ;
      RECT 2.5590 0.7000 2.6090 1.2660 ;
      RECT 2.5590 0.5920 2.6090 0.6500 ;
      RECT 2.2550 0.5420 2.6090 0.5920 ;
      RECT 2.5590 0.3690 2.6090 0.5420 ;
      RECT 1.6310 0.5180 1.7370 0.5680 ;
      RECT 1.6870 0.5680 1.7370 0.6180 ;
      RECT 1.6870 0.6180 2.0930 0.6680 ;
      RECT 1.6870 0.6680 1.7370 0.7510 ;
      RECT 1.6470 0.7510 1.7370 0.8010 ;
      RECT 1.6470 0.8010 1.6970 0.9920 ;
      RECT 1.0390 1.2040 1.2410 1.2540 ;
      RECT 1.0390 0.7500 1.0890 1.2040 ;
      RECT 1.1910 0.5680 1.2410 1.2040 ;
      RECT 1.0390 0.1960 1.0890 0.5180 ;
      RECT 1.1910 0.2820 1.2410 0.5180 ;
      RECT 1.0390 0.5180 1.2410 0.5680 ;
      RECT 3.0550 0.6040 4.3730 0.6540 ;
      RECT 3.0550 0.6540 3.1050 0.8860 ;
      RECT 3.0550 0.5880 3.1050 0.6040 ;
      RECT 3.0150 0.8860 3.1050 0.9360 ;
      RECT 3.0150 0.5630 3.1050 0.5880 ;
      RECT 3.0150 0.9360 3.0650 1.3580 ;
      RECT 3.0150 0.5110 3.1050 0.5130 ;
      RECT 3.0150 0.2820 3.0650 0.5110 ;
      RECT 2.6940 0.5130 3.1050 0.5630 ;
      RECT 0.6430 1.5260 1.6570 1.5760 ;
      RECT 1.6070 1.0920 1.6570 1.5260 ;
      RECT 1.6070 1.0420 1.9250 1.0920 ;
      RECT 1.8750 0.7180 1.9250 1.0420 ;
      RECT 0.2790 0.6180 0.7250 0.6680 ;
      RECT 0.2790 0.6680 0.3290 0.9140 ;
      RECT 0.2790 0.4220 0.3290 0.6180 ;
      RECT 0.7350 0.5180 0.8610 0.5680 ;
      RECT 0.8110 0.5680 0.8610 0.7180 ;
      RECT 0.7350 0.7180 0.8610 0.7680 ;
      RECT 0.7350 0.3940 0.7850 0.5180 ;
      RECT 0.7350 0.7680 0.7850 0.9140 ;
      RECT 2.1430 0.4680 2.1930 0.7280 ;
      RECT 1.9750 0.7280 2.1930 0.7780 ;
      RECT 1.3430 0.6180 1.6370 0.6680 ;
      RECT 1.9750 0.7780 2.0250 1.2200 ;
      RECT 1.7830 1.2200 2.0250 1.2700 ;
      RECT 1.3430 0.4180 2.1930 0.4680 ;
      RECT 1.3430 0.4680 1.3930 0.6180 ;
      RECT 1.3430 0.2820 1.3930 0.4180 ;
      RECT 1.3430 0.6680 1.3930 1.2540 ;
      RECT 1.7070 1.5310 1.9450 1.5810 ;
      RECT 2.0110 1.5310 2.5490 1.5810 ;
      RECT 0.6430 0.0960 2.8530 0.1460 ;
    LAYER PO ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 1.2770 0.9900 1.3070 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 4.6210 0.0680 4.6510 1.6060 ;
      RECT 4.3170 0.0680 4.3470 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 4.4690 0.0680 4.4990 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 1.8850 0.0680 1.9150 0.8120 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 2.0370 0.0680 2.0670 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 1.8850 1.0820 1.9150 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 3.7090 0.0680 3.7390 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 1.2770 0.0680 1.3070 0.6420 ;
  END
END CGLNPSX8_LVT

MACRO CGLPPRX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.496 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 0.0890 0.8770 0.2070 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 3.4960 0.0300 ;
        RECT 2.8230 0.0300 2.8730 0.1970 ;
        RECT 0.2790 0.0300 0.3290 0.3370 ;
        RECT 0.5830 0.0300 0.6330 0.2820 ;
        RECT 3.2090 0.0300 3.2590 0.1970 ;
        RECT 2.2530 0.0300 2.3030 0.1470 ;
        RECT 2.8230 0.1970 2.9130 0.2470 ;
        RECT 0.5830 0.2820 1.0890 0.3320 ;
        RECT 3.1670 0.1970 3.2590 0.2470 ;
        RECT 2.0750 0.1470 2.3030 0.1880 ;
        RECT 2.8630 0.2470 2.9130 0.3710 ;
        RECT 1.0390 0.3320 1.0890 0.5780 ;
        RECT 0.8870 0.3320 0.9370 0.5640 ;
        RECT 1.0390 0.2700 1.0890 0.2820 ;
        RECT 3.1670 0.2470 3.2170 0.3710 ;
        RECT 2.0750 0.1880 2.4730 0.1970 ;
        RECT 1.0390 0.2200 1.6970 0.2700 ;
        RECT 2.2530 0.1970 2.4730 0.2380 ;
        RECT 1.6470 0.2700 1.6970 0.4080 ;
        RECT 1.6470 0.2190 1.6970 0.2200 ;
    END
  END VSS

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4910 0.6130 0.6630 0.6630 ;
        RECT 0.5530 0.5530 0.6630 0.6130 ;
    END
    ANTENNAGATEAREA 0.018 ;
  END SE

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 3.4960 1.7020 ;
        RECT 2.8630 0.9260 2.9130 1.6420 ;
        RECT 3.1670 0.9260 3.2170 1.6420 ;
        RECT 1.3840 1.4560 1.4340 1.6420 ;
        RECT 2.5990 1.2540 2.6490 1.6420 ;
        RECT 0.5830 1.4060 1.4340 1.4560 ;
        RECT 1.6470 1.2040 2.6490 1.2540 ;
        RECT 1.0390 0.7990 1.0890 1.4060 ;
        RECT 0.8870 0.8120 0.9370 1.4060 ;
        RECT 0.5830 0.8060 0.6330 1.4060 ;
        RECT 2.1030 0.7580 2.1530 1.2040 ;
        RECT 2.5590 0.8980 2.6090 1.2040 ;
        RECT 1.6470 0.9000 1.6970 1.2040 ;
    END
  END VDD

  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9850 0.8340 3.1330 0.8840 ;
        RECT 2.9850 0.8840 3.0950 0.9670 ;
        RECT 3.0830 0.4670 3.1330 0.8340 ;
        RECT 3.0150 0.9670 3.0650 1.5610 ;
        RECT 3.0150 0.4170 3.1330 0.4670 ;
        RECT 3.0150 0.1970 3.0650 0.4170 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END GCLK

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2480 1.3130 0.3590 1.3170 ;
        RECT 0.2480 1.3170 0.4210 1.3670 ;
        RECT 0.2480 1.3670 0.3590 1.4230 ;
    END
    ANTENNAGATEAREA 0.018 ;
  END EN
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 3.6110 1.7870 ;
    LAYER M1 ;
      RECT 2.2950 0.6390 2.6850 0.6890 ;
      RECT 2.6350 0.5880 2.6850 0.6390 ;
      RECT 1.7570 0.1380 1.8070 0.3580 ;
      RECT 1.7070 0.0880 1.8070 0.1380 ;
      RECT 2.2950 0.6890 2.3450 0.7550 ;
      RECT 2.2950 0.5510 2.3450 0.6390 ;
      RECT 2.2550 0.7550 2.3450 0.8050 ;
      RECT 2.0510 0.5010 2.3450 0.5510 ;
      RECT 2.2550 0.8050 2.3050 1.1130 ;
      RECT 2.2550 0.4690 2.3050 0.5010 ;
      RECT 2.0510 0.4080 2.1010 0.5010 ;
      RECT 1.7570 0.3580 2.1010 0.4080 ;
      RECT 0.7350 0.6640 1.0290 0.7140 ;
      RECT 0.7350 0.7140 0.7850 1.2310 ;
      RECT 0.7350 0.4500 0.7850 0.6640 ;
      RECT 1.9510 0.6350 2.2450 0.6850 ;
      RECT 1.4940 0.5090 1.5440 0.5170 ;
      RECT 1.4940 0.3630 1.5440 0.4590 ;
      RECT 1.4430 0.5170 1.5440 0.5670 ;
      RECT 1.4430 0.5670 1.4930 0.8340 ;
      RECT 1.4430 0.8340 1.5440 0.8840 ;
      RECT 1.4940 0.8840 1.5440 1.1600 ;
      RECT 1.9510 0.5090 2.0010 0.6350 ;
      RECT 1.9910 0.6850 2.0410 0.8360 ;
      RECT 1.4940 0.4590 2.0010 0.5090 ;
      RECT 1.9510 0.8360 2.0410 0.8860 ;
      RECT 1.9510 0.4580 2.0010 0.4590 ;
      RECT 1.9510 0.8860 2.0010 1.1120 ;
      RECT 2.7960 0.6610 3.0050 0.7110 ;
      RECT 2.7960 0.7110 2.8460 0.7560 ;
      RECT 2.7960 0.5380 2.8460 0.6610 ;
      RECT 2.4070 0.7560 2.8460 0.8060 ;
      RECT 2.7110 0.4880 2.8460 0.5380 ;
      RECT 2.4070 0.8060 2.4570 1.1140 ;
      RECT 2.7110 0.8060 2.7610 1.1140 ;
      RECT 2.7110 0.1900 2.7610 0.4880 ;
      RECT 1.5360 1.5340 2.5490 1.5840 ;
      RECT 1.1910 0.8500 1.2410 1.2500 ;
      RECT 1.1470 0.8000 1.2410 0.8500 ;
      RECT 1.1470 0.5940 1.1970 0.8000 ;
      RECT 1.1470 0.5440 1.2410 0.5940 ;
      RECT 1.1910 0.3280 1.2410 0.5440 ;
      RECT 1.5360 1.3000 1.5860 1.5340 ;
      RECT 1.1910 1.2500 1.5860 1.3000 ;
      RECT 0.4710 1.5260 1.3330 1.5760 ;
      RECT 0.2790 1.1870 0.5210 1.2370 ;
      RECT 0.2790 0.5030 0.3290 1.1870 ;
      RECT 0.2790 0.4530 0.4810 0.5030 ;
      RECT 0.4310 0.2370 0.4810 0.4530 ;
      RECT 0.4710 1.2370 0.5210 1.5260 ;
      RECT 0.9470 0.0950 1.6370 0.1450 ;
      RECT 2.9230 0.0970 3.1580 0.1470 ;
      RECT 2.1550 0.3690 2.6340 0.4190 ;
      RECT 2.5840 0.1380 2.6340 0.3690 ;
      RECT 2.1550 0.3080 2.2050 0.3690 ;
      RECT 2.4610 0.0880 2.6340 0.1380 ;
      RECT 1.8750 0.2880 2.2050 0.3080 ;
      RECT 1.8750 0.2580 2.2030 0.2880 ;
      RECT 1.8750 0.0880 1.9250 0.2580 ;
      RECT 1.3430 0.6950 1.3930 1.1240 ;
      RECT 1.2470 0.6450 1.3930 0.6950 ;
      RECT 1.3430 0.3630 1.3930 0.6450 ;
      RECT 1.5710 0.7850 1.6210 0.7870 ;
      RECT 1.5710 0.7350 1.9410 0.7850 ;
      RECT 1.5710 0.6270 1.6210 0.7350 ;
    LAYER PO ;
      RECT 1.2770 0.0840 1.3070 1.6060 ;
      RECT 0.6690 0.0900 0.6990 1.6060 ;
      RECT 1.4290 0.6900 1.4590 1.5900 ;
      RECT 1.5810 0.0880 1.6110 1.5900 ;
      RECT 0.2130 0.1100 0.2430 1.6060 ;
      RECT 0.3650 0.1080 0.3950 1.6060 ;
      RECT 0.0610 0.1100 0.0910 1.6060 ;
      RECT 2.7970 0.0670 2.8270 1.6080 ;
      RECT 3.1010 0.0860 3.1310 1.6100 ;
      RECT 1.7330 0.0780 1.7630 1.5900 ;
      RECT 1.8850 0.6900 1.9150 1.5900 ;
      RECT 1.4290 0.0850 1.4590 0.5900 ;
      RECT 1.8850 0.0780 1.9150 0.5900 ;
      RECT 2.9490 0.0860 2.9790 1.6100 ;
      RECT 3.2530 0.0880 3.2830 1.5900 ;
      RECT 2.4930 0.0760 2.5230 1.6060 ;
      RECT 3.4050 0.0880 3.4350 1.5900 ;
      RECT 2.1890 0.0810 2.2190 1.5900 ;
      RECT 2.6450 0.0760 2.6750 1.6060 ;
      RECT 2.0370 0.0810 2.0670 1.5900 ;
      RECT 0.5170 0.1080 0.5470 1.6060 ;
      RECT 2.3410 0.0810 2.3710 1.5900 ;
      RECT 1.1250 0.0840 1.1550 1.6060 ;
      RECT 0.9730 0.0840 1.0030 1.6060 ;
      RECT 0.8210 0.0840 0.8510 1.6060 ;
  END
END CGLPPRX2_LVT

MACRO CGLPPRX8_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.408 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2480 1.3130 0.3590 1.3170 ;
        RECT 0.2480 1.3170 0.4210 1.3670 ;
        RECT 0.2480 1.3670 0.3590 1.4230 ;
    END
    ANTENNAGATEAREA 0.018 ;
  END EN

  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9850 0.8340 3.1330 0.8840 ;
        RECT 2.9850 0.8840 3.0950 0.9670 ;
        RECT 3.0830 0.7030 3.1330 0.8340 ;
        RECT 3.0150 0.9670 3.0650 1.5610 ;
        RECT 3.0830 0.6530 3.9770 0.7030 ;
        RECT 3.0830 0.5790 3.1330 0.6530 ;
        RECT 3.9270 0.7030 3.9770 1.5700 ;
        RECT 3.9270 0.3480 3.9770 0.6530 ;
        RECT 3.6230 0.7030 3.6730 1.5600 ;
        RECT 3.6230 0.3480 3.6730 0.6530 ;
        RECT 3.3190 0.7030 3.3690 1.5600 ;
        RECT 3.3190 0.3480 3.3690 0.6530 ;
        RECT 3.0150 0.5290 3.1330 0.5790 ;
        RECT 3.0150 0.3130 3.0650 0.5290 ;
    END
    ANTENNADIFFAREA 0.5952 ;
  END GCLK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.4080 1.7020 ;
        RECT 3.1670 0.9260 3.2170 1.6420 ;
        RECT 4.0790 0.8340 4.1290 1.6420 ;
        RECT 3.7750 0.8340 3.8250 1.6420 ;
        RECT 3.4710 0.8340 3.5210 1.6420 ;
        RECT 2.8630 0.9260 2.9130 1.6420 ;
        RECT 1.3840 1.4560 1.4340 1.6420 ;
        RECT 2.5990 1.2540 2.6490 1.6420 ;
        RECT 0.5830 1.4060 1.4340 1.4560 ;
        RECT 1.6470 1.2040 2.6490 1.2540 ;
        RECT 1.0390 0.7990 1.0890 1.4060 ;
        RECT 0.5830 0.8100 0.6330 1.4060 ;
        RECT 0.8870 0.8120 0.9370 1.4060 ;
        RECT 2.1030 0.7580 2.1530 1.2040 ;
        RECT 2.5590 0.8980 2.6090 1.2040 ;
        RECT 1.6470 0.9000 1.6970 1.2040 ;
    END
  END VDD

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4910 0.6130 0.6630 0.6630 ;
        RECT 0.5530 0.5530 0.6630 0.6130 ;
    END
    ANTENNAGATEAREA 0.018 ;
  END SE

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.4080 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.3370 ;
        RECT 0.5830 0.0300 0.6330 0.2820 ;
        RECT 2.8230 0.0300 2.8730 0.1970 ;
        RECT 2.2530 0.0300 2.3030 0.1470 ;
        RECT 0.5830 0.2820 1.0890 0.3320 ;
        RECT 2.8230 0.1970 4.1290 0.2470 ;
        RECT 2.0750 0.1470 2.3030 0.1890 ;
        RECT 0.8870 0.3320 0.9370 0.5320 ;
        RECT 1.0390 0.3320 1.0890 0.5460 ;
        RECT 1.0390 0.2380 1.0890 0.2820 ;
        RECT 3.1670 0.2470 3.2170 0.3710 ;
        RECT 4.0790 0.2470 4.1290 0.5610 ;
        RECT 3.4710 0.2470 3.5210 0.5610 ;
        RECT 3.7750 0.2470 3.8250 0.5610 ;
        RECT 2.8630 0.2470 2.9130 0.3710 ;
        RECT 2.0750 0.1890 2.4730 0.1970 ;
        RECT 1.0390 0.1880 1.6970 0.2380 ;
        RECT 2.2530 0.1970 2.4730 0.2390 ;
        RECT 1.6470 0.2380 1.6970 0.4080 ;
    END
  END VSS

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 0.0960 0.8770 0.2250 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 4.5230 1.7870 ;
    LAYER M1 ;
      RECT 2.2950 0.6390 2.6850 0.6890 ;
      RECT 2.6350 0.5880 2.6850 0.6390 ;
      RECT 2.2950 0.6890 2.3450 0.7550 ;
      RECT 2.2950 0.5510 2.3450 0.6390 ;
      RECT 2.2550 0.7550 2.3450 0.8050 ;
      RECT 2.0510 0.5010 2.3450 0.5510 ;
      RECT 2.2550 0.8050 2.3050 1.1130 ;
      RECT 2.2550 0.4690 2.3050 0.5010 ;
      RECT 1.7570 0.1380 1.8070 0.3580 ;
      RECT 1.7070 0.0880 1.8070 0.1380 ;
      RECT 2.0510 0.4080 2.1010 0.5010 ;
      RECT 1.7570 0.3580 2.1010 0.4080 ;
      RECT 2.1550 0.3690 2.6340 0.4190 ;
      RECT 2.5840 0.1390 2.6340 0.3690 ;
      RECT 2.1550 0.3080 2.2050 0.3690 ;
      RECT 2.4620 0.0890 2.6350 0.1390 ;
      RECT 1.8750 0.2890 2.2050 0.3080 ;
      RECT 1.8750 0.2580 2.2030 0.2890 ;
      RECT 1.8750 0.0880 1.9250 0.2580 ;
      RECT 2.7960 0.6610 3.0050 0.7110 ;
      RECT 2.7960 0.5380 2.8460 0.6610 ;
      RECT 2.7960 0.7110 2.8460 0.7560 ;
      RECT 2.6950 0.4880 2.8460 0.5380 ;
      RECT 2.4070 0.7560 2.8460 0.8060 ;
      RECT 2.4070 0.8060 2.4570 1.0220 ;
      RECT 2.7110 0.1910 2.7610 0.4880 ;
      RECT 2.7110 0.8060 2.7610 1.0220 ;
      RECT 0.4710 1.5260 1.3330 1.5760 ;
      RECT 0.2790 1.1870 0.5210 1.2370 ;
      RECT 0.4710 1.2370 0.5210 1.5260 ;
      RECT 0.2790 0.5030 0.3290 1.1870 ;
      RECT 0.2790 0.4530 0.4810 0.5030 ;
      RECT 0.4310 0.2370 0.4810 0.4530 ;
      RECT 1.5360 1.5340 2.5490 1.5840 ;
      RECT 1.1910 0.8500 1.2410 1.2500 ;
      RECT 1.1470 0.8000 1.2410 0.8500 ;
      RECT 1.1470 0.5680 1.1970 0.8000 ;
      RECT 1.1470 0.5180 1.2410 0.5680 ;
      RECT 1.1910 0.3020 1.2410 0.5180 ;
      RECT 1.5360 1.3000 1.5860 1.5340 ;
      RECT 1.1910 1.2500 1.5860 1.3000 ;
      RECT 1.5360 1.2480 1.5860 1.2500 ;
      RECT 2.9230 0.0970 4.0690 0.1470 ;
      RECT 1.9510 0.6350 2.2450 0.6850 ;
      RECT 1.9510 0.5090 2.0010 0.6350 ;
      RECT 1.9910 0.6850 2.0410 0.8360 ;
      RECT 1.4940 0.4590 2.0010 0.5090 ;
      RECT 1.9510 0.8360 2.0410 0.8860 ;
      RECT 1.9510 0.4580 2.0010 0.4590 ;
      RECT 1.9510 0.8860 2.0010 1.1120 ;
      RECT 1.4940 0.5090 1.5440 0.5170 ;
      RECT 1.4940 0.3630 1.5440 0.4590 ;
      RECT 1.4430 0.5170 1.5440 0.5670 ;
      RECT 1.4430 0.5670 1.4930 0.8340 ;
      RECT 1.4430 0.8340 1.5440 0.8840 ;
      RECT 1.4940 0.8840 1.5440 1.1600 ;
      RECT 0.9470 0.0880 1.6370 0.1380 ;
      RECT 0.7350 0.6180 1.0290 0.6680 ;
      RECT 0.7350 0.6680 0.7850 1.1900 ;
      RECT 0.7350 0.4180 0.7850 0.6180 ;
      RECT 1.2470 0.6450 1.3930 0.6950 ;
      RECT 1.3430 0.6950 1.3930 1.1240 ;
      RECT 1.3430 0.3630 1.3930 0.6450 ;
      RECT 1.5710 0.7350 1.9410 0.7850 ;
      RECT 1.5710 0.7850 1.6210 0.7870 ;
      RECT 1.5710 0.6270 1.6210 0.7350 ;
    LAYER PO ;
      RECT 3.2530 0.0860 3.2830 1.6100 ;
      RECT 2.7970 0.0940 2.8270 1.6080 ;
      RECT 0.0610 0.1100 0.0910 1.6060 ;
      RECT 0.3650 0.1080 0.3950 1.6060 ;
      RECT 0.2130 0.1100 0.2430 1.6060 ;
      RECT 1.5810 0.0740 1.6110 1.5900 ;
      RECT 1.4290 0.6900 1.4590 1.5900 ;
      RECT 0.6690 0.0660 0.6990 1.6060 ;
      RECT 1.2770 0.0680 1.3070 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 2.3410 0.0810 2.3710 1.5900 ;
      RECT 0.5170 0.1080 0.5470 1.6060 ;
      RECT 2.0370 0.0810 2.0670 1.5900 ;
      RECT 2.6450 0.1190 2.6750 1.6060 ;
      RECT 2.1890 0.0810 2.2190 1.5900 ;
      RECT 4.3170 0.1020 4.3470 1.5900 ;
      RECT 2.4930 0.0710 2.5230 1.6060 ;
      RECT 4.1650 0.1020 4.1950 1.5900 ;
      RECT 2.9490 0.0860 2.9790 1.6100 ;
      RECT 1.8850 0.0740 1.9150 0.5900 ;
      RECT 1.4290 0.0710 1.4590 0.5900 ;
      RECT 1.8850 0.6900 1.9150 1.5900 ;
      RECT 1.7330 0.0740 1.7630 1.5900 ;
      RECT 3.1010 0.0860 3.1310 1.6100 ;
      RECT 3.8610 0.0860 3.8910 1.6100 ;
      RECT 4.0130 0.0860 4.0430 1.6100 ;
      RECT 3.4050 0.0860 3.4350 1.6100 ;
      RECT 3.5570 0.0860 3.5870 1.6100 ;
      RECT 3.7090 0.0860 3.7390 1.6100 ;
  END
END CGLPPRX8_LVT

MACRO CGLPPSX16_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.232 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.5990 0.1480 5.6490 0.5040 ;
        RECT 3.4710 0.5040 6.0350 0.5530 ;
        RECT 5.9030 0.1480 5.9530 0.5040 ;
        RECT 5.2950 0.1480 5.3450 0.5040 ;
        RECT 4.9910 0.1480 5.0410 0.5040 ;
        RECT 4.6870 0.1480 4.7370 0.5040 ;
        RECT 4.3830 0.1480 4.4330 0.5040 ;
        RECT 4.0790 0.1480 4.1290 0.5040 ;
        RECT 3.7750 0.1480 3.8250 0.5040 ;
        RECT 3.4710 0.1480 3.5210 0.5040 ;
        RECT 3.4710 0.5530 6.1350 0.5540 ;
        RECT 5.9850 0.5540 6.1350 0.6630 ;
        RECT 5.9850 0.6630 6.0350 0.8040 ;
        RECT 3.4710 0.8040 6.0350 0.8540 ;
        RECT 5.5990 0.8540 5.6490 1.5460 ;
        RECT 5.9030 0.8540 5.9530 1.5460 ;
        RECT 5.2950 0.8540 5.3450 1.5460 ;
        RECT 4.9910 0.8540 5.0410 1.5460 ;
        RECT 4.6870 0.8540 4.7370 1.5460 ;
        RECT 4.3830 0.8540 4.4330 1.5460 ;
        RECT 4.0790 0.8540 4.1290 1.5460 ;
        RECT 3.7750 0.8540 3.8250 1.5460 ;
        RECT 3.4710 0.8540 3.5210 1.5460 ;
    END
    ANTENNADIFFAREA 1.2904 ;
  END GCLK

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 0.8570 0.9670 0.9670 ;
        RECT 0.9170 0.6680 0.9670 0.8570 ;
        RECT 0.9170 0.6180 1.0290 0.6680 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END EN

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2250 0.6180 2.3970 0.6680 ;
        RECT 2.2250 0.5530 2.3350 0.6180 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END SE

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 6.2320 1.7020 ;
        RECT 3.9270 0.9040 3.9770 1.6420 ;
        RECT 3.6230 0.9040 3.6730 1.6420 ;
        RECT 4.2310 0.9040 4.2810 1.6420 ;
        RECT 5.7510 0.9040 5.8010 1.6420 ;
        RECT 5.1430 0.9040 5.1930 1.6420 ;
        RECT 4.8390 0.9040 4.8890 1.6420 ;
        RECT 5.4470 0.9040 5.4970 1.6420 ;
        RECT 4.5350 0.9040 4.5850 1.6420 ;
        RECT 0.5830 1.3540 0.6330 1.6420 ;
        RECT 3.1670 1.3660 3.2170 1.6420 ;
        RECT 2.2710 1.3850 2.3210 1.6420 ;
        RECT 0.4310 1.3040 1.5450 1.3540 ;
        RECT 2.6950 1.3160 3.2170 1.3660 ;
        RECT 1.7990 1.3350 2.3210 1.3850 ;
        RECT 0.4310 1.0880 0.4810 1.3040 ;
        RECT 1.4950 0.7500 1.5450 1.3040 ;
        RECT 0.8870 1.0370 0.9370 1.3040 ;
        RECT 0.5830 1.1010 0.6330 1.3040 ;
        RECT 3.1670 1.2660 3.2170 1.3160 ;
        RECT 1.7990 1.1420 1.8490 1.3350 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 6.2320 0.0300 ;
        RECT 3.6230 0.0300 3.6730 0.4540 ;
        RECT 3.9270 0.0300 3.9770 0.4540 ;
        RECT 4.2310 0.0300 4.2810 0.4540 ;
        RECT 4.5350 0.0300 4.5850 0.4540 ;
        RECT 4.8390 0.0300 4.8890 0.4540 ;
        RECT 5.1430 0.0300 5.1930 0.4540 ;
        RECT 5.4470 0.0300 5.4970 0.4540 ;
        RECT 5.7510 0.0300 5.8010 0.4540 ;
        RECT 0.4310 0.0300 0.4810 0.1960 ;
        RECT 1.8390 0.0300 1.8890 0.3180 ;
        RECT 0.4310 0.1960 0.9370 0.2460 ;
        RECT 1.4790 0.3180 2.3050 0.3680 ;
        RECT 0.4310 0.2460 0.4810 0.4500 ;
        RECT 0.5830 0.2460 0.6330 0.4500 ;
        RECT 0.8870 0.2460 0.9370 0.4500 ;
        RECT 2.2550 0.3680 2.3050 0.4830 ;
        RECT 2.2550 0.2460 2.3050 0.3180 ;
        RECT 2.2550 0.1960 3.0650 0.2460 ;
        RECT 3.0150 0.2460 3.0650 0.5820 ;
        RECT 2.5590 0.2460 2.6090 0.4680 ;
    END
  END VSS

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 1.4240 0.4210 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 6.3470 1.7870 ;
    LAYER M1 ;
      RECT 2.0110 0.0960 3.1570 0.1460 ;
      RECT 0.2790 0.6180 0.7250 0.6680 ;
      RECT 0.2790 0.6680 0.3290 0.9140 ;
      RECT 0.2790 0.4220 0.3290 0.6180 ;
      RECT 0.6430 0.0960 1.7890 0.1460 ;
      RECT 2.8630 0.7860 3.3090 0.8360 ;
      RECT 2.9030 0.5680 2.9530 0.7860 ;
      RECT 2.8630 0.8360 2.9130 1.1030 ;
      RECT 2.8630 0.5180 2.9530 0.5680 ;
      RECT 2.5420 1.1030 2.9130 1.1530 ;
      RECT 2.8630 0.2960 2.9130 0.5180 ;
      RECT 2.8630 1.1530 2.9130 1.2660 ;
      RECT 1.6470 0.7510 1.7370 0.8010 ;
      RECT 1.6470 0.8010 1.6970 0.9920 ;
      RECT 1.6870 0.6680 1.7370 0.7510 ;
      RECT 1.6870 0.6180 1.9410 0.6680 ;
      RECT 1.6870 0.5680 1.7370 0.6180 ;
      RECT 1.6310 0.5180 1.7370 0.5680 ;
      RECT 0.7350 0.5180 0.8610 0.5680 ;
      RECT 0.8110 0.5680 0.8610 0.7180 ;
      RECT 0.7350 0.7180 0.8610 0.7680 ;
      RECT 0.7350 0.3940 0.7850 0.5180 ;
      RECT 0.7350 0.7680 0.7850 0.9140 ;
      RECT 2.4940 0.6180 2.8530 0.6680 ;
      RECT 2.4940 0.6680 2.5440 0.7200 ;
      RECT 2.4940 0.5680 2.5440 0.6180 ;
      RECT 2.4070 0.7200 2.5440 0.7700 ;
      RECT 2.4070 0.5180 2.5440 0.5680 ;
      RECT 2.4070 0.7700 2.4570 1.1620 ;
      RECT 2.4070 0.3940 2.4570 0.5180 ;
      RECT 3.3190 0.6040 5.8930 0.6540 ;
      RECT 3.3190 0.2820 3.3690 0.6040 ;
      RECT 3.3590 0.6540 3.4090 0.8860 ;
      RECT 3.3190 0.8860 3.4090 0.9360 ;
      RECT 3.3190 0.9360 3.3690 1.1660 ;
      RECT 3.3190 1.2160 3.3690 1.3580 ;
      RECT 2.9980 1.1660 3.3690 1.2160 ;
      RECT 2.5620 1.4280 2.7010 1.4780 ;
      RECT 2.5620 1.2700 2.6120 1.4280 ;
      RECT 2.0870 1.2200 2.6120 1.2700 ;
      RECT 1.3430 0.2820 1.3930 0.4180 ;
      RECT 1.3430 0.4680 1.3930 0.6180 ;
      RECT 1.3430 0.6680 1.3930 1.2540 ;
      RECT 1.3430 0.6180 1.6370 0.6680 ;
      RECT 2.1030 0.4680 2.1530 0.7280 ;
      RECT 1.3430 0.4180 2.1530 0.4680 ;
      RECT 2.2380 0.7780 2.2880 1.2200 ;
      RECT 2.1030 0.7280 2.2880 0.7780 ;
      RECT 1.9760 0.8280 2.0930 0.8780 ;
      RECT 1.9760 0.8780 2.0260 1.0420 ;
      RECT 1.6070 1.0420 2.0260 1.0920 ;
      RECT 1.6070 1.0920 1.6570 1.5260 ;
      RECT 0.7950 1.5260 1.6570 1.5760 ;
      RECT 1.0390 0.1960 1.0890 0.5180 ;
      RECT 1.1910 0.2820 1.2410 0.5180 ;
      RECT 1.1910 0.5680 1.2410 1.2040 ;
      RECT 1.0390 1.2040 1.2410 1.2540 ;
      RECT 1.0390 0.7500 1.0890 1.2040 ;
      RECT 1.0390 0.5180 1.2410 0.5680 ;
      RECT 1.7070 1.5310 2.0930 1.5810 ;
    LAYER PO ;
      RECT 2.0370 0.0680 2.0670 0.9060 ;
      RECT 5.9890 0.0680 6.0190 1.6060 ;
      RECT 5.8370 0.0680 5.8670 1.6060 ;
      RECT 5.0770 0.0680 5.1070 1.6060 ;
      RECT 4.9250 0.0680 4.9550 1.6060 ;
      RECT 4.7730 0.0680 4.8030 1.6060 ;
      RECT 4.6210 0.0680 4.6510 1.6060 ;
      RECT 5.3810 0.0680 5.4110 1.6060 ;
      RECT 5.2290 0.0680 5.2590 1.6060 ;
      RECT 5.5330 0.0680 5.5630 1.6060 ;
      RECT 4.4690 0.0680 4.4990 1.6060 ;
      RECT 4.3170 0.0680 4.3470 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 2.0370 1.0820 2.0670 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 3.7090 0.0680 3.7390 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 6.1410 0.0680 6.1710 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 1.2770 0.0680 1.3070 0.6420 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 1.2770 0.9900 1.3070 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 5.6850 0.0680 5.7150 1.6060 ;
  END
END CGLPPSX16_LVT

MACRO CGLPPSX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.104 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 0.8570 0.9670 0.9670 ;
        RECT 0.9170 0.6680 0.9670 0.8570 ;
        RECT 0.9170 0.6180 1.0290 0.6680 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END EN

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2250 0.5530 2.3350 0.6180 ;
        RECT 2.2250 0.6180 2.3970 0.6680 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END SE

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.1040 1.7020 ;
        RECT 3.6230 0.9040 3.6730 1.6420 ;
        RECT 0.5830 1.3540 0.6330 1.6420 ;
        RECT 3.1670 1.3660 3.2170 1.6420 ;
        RECT 2.2710 1.3850 2.3210 1.6420 ;
        RECT 0.4310 1.3040 1.5450 1.3540 ;
        RECT 2.6950 1.3160 3.2170 1.3660 ;
        RECT 1.7990 1.3350 2.3210 1.3850 ;
        RECT 0.4310 1.0880 0.4810 1.3040 ;
        RECT 1.4950 0.7500 1.5450 1.3040 ;
        RECT 0.8870 1.0370 0.9370 1.3040 ;
        RECT 0.5830 1.1010 0.6330 1.3040 ;
        RECT 3.1670 1.2660 3.2170 1.3160 ;
        RECT 1.7990 1.1420 1.8490 1.3350 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.1040 0.0300 ;
        RECT 3.6230 0.0300 3.6730 0.4540 ;
        RECT 0.4310 0.0300 0.4810 0.1960 ;
        RECT 1.8390 0.0300 1.8890 0.3180 ;
        RECT 0.4310 0.1960 0.9370 0.2460 ;
        RECT 1.4790 0.3180 2.3050 0.3680 ;
        RECT 0.4310 0.2460 0.4810 0.4500 ;
        RECT 0.8870 0.2460 0.9370 0.4500 ;
        RECT 0.5830 0.2460 0.6330 0.4500 ;
        RECT 2.2550 0.3680 2.3050 0.4830 ;
        RECT 2.2550 0.2460 2.3050 0.3180 ;
        RECT 2.2550 0.1960 3.0650 0.2460 ;
        RECT 2.5590 0.2460 2.6090 0.4080 ;
        RECT 3.0150 0.2460 3.0650 0.5820 ;
    END
  END VSS

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 1.4240 0.4210 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.7450 1.0090 3.8650 1.1190 ;
        RECT 3.7750 1.1190 3.8250 1.5460 ;
        RECT 3.8150 0.8540 3.8650 1.0090 ;
        RECT 3.4710 0.8040 3.8650 0.8540 ;
        RECT 3.4710 0.8540 3.5210 1.5460 ;
        RECT 3.8150 0.5540 3.8650 0.8040 ;
        RECT 3.4710 0.5040 3.8650 0.5540 ;
        RECT 3.7750 0.1480 3.8250 0.5040 ;
        RECT 3.4710 0.1480 3.5210 0.5040 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END GCLK
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 4.2190 1.7870 ;
    LAYER M1 ;
      RECT 2.8630 0.7860 3.3090 0.8360 ;
      RECT 2.9030 0.5020 2.9530 0.7860 ;
      RECT 2.8630 0.8360 2.9130 1.1030 ;
      RECT 2.8630 0.4520 2.9530 0.5020 ;
      RECT 2.5420 1.1030 2.9130 1.1530 ;
      RECT 2.8630 0.3130 2.9130 0.4520 ;
      RECT 2.8630 1.1530 2.9130 1.2660 ;
      RECT 3.3190 0.6040 3.7650 0.6540 ;
      RECT 3.3190 0.2820 3.3690 0.6040 ;
      RECT 3.3590 0.6540 3.4090 0.8860 ;
      RECT 3.3190 0.8860 3.4090 0.9360 ;
      RECT 3.3190 0.9360 3.3690 1.1660 ;
      RECT 3.3190 1.2160 3.3690 1.3580 ;
      RECT 2.9980 1.1660 3.3690 1.2160 ;
      RECT 0.2790 0.6180 0.7250 0.6680 ;
      RECT 0.2790 0.6680 0.3290 0.9140 ;
      RECT 0.2790 0.4220 0.3290 0.6180 ;
      RECT 0.7350 0.5180 0.8610 0.5680 ;
      RECT 0.8110 0.5680 0.8610 0.7180 ;
      RECT 0.7350 0.7180 0.8610 0.7680 ;
      RECT 0.7350 0.3940 0.7850 0.5180 ;
      RECT 0.7350 0.7680 0.7850 0.9140 ;
      RECT 1.6470 0.7510 1.7370 0.8010 ;
      RECT 1.6470 0.8010 1.6970 0.9920 ;
      RECT 1.6870 0.6680 1.7370 0.7510 ;
      RECT 1.6870 0.6180 1.9410 0.6680 ;
      RECT 1.6870 0.5680 1.7370 0.6180 ;
      RECT 1.6310 0.5180 1.7370 0.5680 ;
      RECT 2.5620 1.4280 2.7010 1.4780 ;
      RECT 2.5620 1.2700 2.6120 1.4280 ;
      RECT 2.0870 1.2200 2.6120 1.2700 ;
      RECT 1.3430 0.4680 1.3930 0.6180 ;
      RECT 1.3430 0.2820 1.3930 0.4180 ;
      RECT 1.3430 0.6680 1.3930 1.2540 ;
      RECT 1.3430 0.6180 1.6370 0.6680 ;
      RECT 2.1030 0.4680 2.1530 0.7280 ;
      RECT 1.3430 0.4180 2.1530 0.4680 ;
      RECT 2.2380 0.7780 2.2880 1.2200 ;
      RECT 2.1030 0.7280 2.2880 0.7780 ;
      RECT 1.0390 1.2040 1.2410 1.2540 ;
      RECT 1.0390 0.7500 1.0890 1.2040 ;
      RECT 1.1910 0.5690 1.2410 1.2040 ;
      RECT 1.1910 0.2820 1.2410 0.5190 ;
      RECT 1.0390 0.1960 1.0890 0.5190 ;
      RECT 1.0390 0.5190 1.2410 0.5680 ;
      RECT 1.0790 0.5680 1.2410 0.5690 ;
      RECT 2.4940 0.6180 2.8530 0.6680 ;
      RECT 2.4940 0.5680 2.5440 0.6180 ;
      RECT 2.4940 0.6680 2.5440 0.7200 ;
      RECT 2.4070 0.7200 2.5440 0.7700 ;
      RECT 2.4070 0.5180 2.5440 0.5680 ;
      RECT 2.4070 0.3940 2.4570 0.5180 ;
      RECT 2.4070 0.7700 2.4570 1.1620 ;
      RECT 1.9760 0.8780 2.0260 1.0420 ;
      RECT 1.9760 0.8280 2.0930 0.8780 ;
      RECT 1.6070 1.0420 2.0260 1.0920 ;
      RECT 1.6070 1.0920 1.6570 1.5260 ;
      RECT 0.7950 1.5260 1.6570 1.5760 ;
      RECT 0.6430 0.0960 1.7890 0.1460 ;
      RECT 1.7070 1.5310 2.0930 1.5810 ;
      RECT 2.0110 0.0960 3.1570 0.1460 ;
    LAYER PO ;
      RECT 1.2770 0.9900 1.3070 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 2.0370 0.0680 2.0670 0.9060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 2.0370 1.0820 2.0670 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 3.7090 0.0680 3.7390 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 1.2770 0.0680 1.3070 0.6420 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
  END
END CGLPPSX2_LVT

MACRO CGLPPSX4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.408 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 0.8570 0.9670 0.9670 ;
        RECT 0.9170 0.6680 0.9670 0.8570 ;
        RECT 0.9170 0.6180 1.0290 0.6680 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END EN

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2250 0.5530 2.3350 0.6180 ;
        RECT 2.2250 0.6180 2.3970 0.6680 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END SE

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 4.4080 1.7020 ;
        RECT 3.9270 0.9040 3.9770 1.6420 ;
        RECT 3.6230 0.9040 3.6730 1.6420 ;
        RECT 0.5830 1.3540 0.6330 1.6420 ;
        RECT 3.1670 1.3660 3.2170 1.6420 ;
        RECT 2.2710 1.3850 2.3210 1.6420 ;
        RECT 0.4310 1.3040 1.5450 1.3540 ;
        RECT 2.6950 1.3160 3.2170 1.3660 ;
        RECT 1.7990 1.3350 2.3210 1.3850 ;
        RECT 0.4310 1.0880 0.4810 1.3040 ;
        RECT 1.4950 0.7500 1.5450 1.3040 ;
        RECT 0.8870 1.0370 0.9370 1.3040 ;
        RECT 0.5830 1.1010 0.6330 1.3040 ;
        RECT 3.1670 1.2660 3.2170 1.3160 ;
        RECT 1.7990 1.1420 1.8490 1.3350 ;
    END
  END VDD

  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.4710 0.8040 4.2110 0.8540 ;
        RECT 4.0790 0.8540 4.1290 1.5460 ;
        RECT 3.7750 0.8540 3.8250 1.5460 ;
        RECT 3.4710 0.8540 3.5210 1.5460 ;
        RECT 4.1610 0.6630 4.2110 0.8040 ;
        RECT 4.1610 0.5540 4.3110 0.6630 ;
        RECT 3.4710 0.5530 4.3110 0.5540 ;
        RECT 3.4710 0.5040 4.2110 0.5530 ;
        RECT 3.7750 0.1480 3.8250 0.5040 ;
        RECT 4.0790 0.1480 4.1290 0.5040 ;
        RECT 3.4710 0.1480 3.5210 0.5040 ;
    END
    ANTENNADIFFAREA 0.3976 ;
  END GCLK

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 4.4080 0.0300 ;
        RECT 3.9270 0.0300 3.9770 0.4540 ;
        RECT 3.6230 0.0300 3.6730 0.4540 ;
        RECT 0.4310 0.0300 0.4810 0.1960 ;
        RECT 1.8390 0.0300 1.8890 0.3180 ;
        RECT 0.4310 0.1960 0.9370 0.2460 ;
        RECT 1.4790 0.3180 2.3050 0.3680 ;
        RECT 0.4310 0.2460 0.4810 0.4500 ;
        RECT 0.8870 0.2460 0.9370 0.4500 ;
        RECT 0.5830 0.2460 0.6330 0.4500 ;
        RECT 2.2550 0.3680 2.3050 0.4830 ;
        RECT 2.2550 0.2460 2.3050 0.3180 ;
        RECT 2.2550 0.1960 3.0650 0.2460 ;
        RECT 2.5590 0.2460 2.6090 0.4680 ;
        RECT 3.0150 0.2460 3.0650 0.5820 ;
    END
  END VSS

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 1.4240 0.4210 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 4.5230 1.7870 ;
    LAYER M1 ;
      RECT 2.8630 0.7860 3.3090 0.8360 ;
      RECT 2.9030 0.5680 2.9530 0.7860 ;
      RECT 2.8630 0.8360 2.9130 1.1030 ;
      RECT 2.8630 0.5180 2.9530 0.5680 ;
      RECT 2.5420 1.1030 2.9130 1.1530 ;
      RECT 2.8630 0.2960 2.9130 0.5180 ;
      RECT 2.8630 1.1530 2.9130 1.2660 ;
      RECT 3.3190 0.6040 4.0690 0.6540 ;
      RECT 3.3190 0.2820 3.3690 0.6040 ;
      RECT 3.3590 0.6540 3.4090 0.8860 ;
      RECT 3.3190 0.8860 3.4090 0.9360 ;
      RECT 3.3190 0.9360 3.3690 1.1660 ;
      RECT 3.3190 1.2160 3.3690 1.3580 ;
      RECT 2.9980 1.1660 3.3690 1.2160 ;
      RECT 2.4940 0.6180 2.8530 0.6680 ;
      RECT 2.4940 0.6680 2.5440 0.7200 ;
      RECT 2.4940 0.5680 2.5440 0.6180 ;
      RECT 2.4070 0.7200 2.5440 0.7700 ;
      RECT 2.4070 0.5180 2.5440 0.5680 ;
      RECT 2.4070 0.7700 2.4570 1.1620 ;
      RECT 2.4070 0.3940 2.4570 0.5180 ;
      RECT 1.9760 0.8780 2.0260 1.0420 ;
      RECT 1.9760 0.8280 2.0930 0.8780 ;
      RECT 1.6070 1.0420 2.0260 1.0920 ;
      RECT 1.6070 1.0920 1.6570 1.5260 ;
      RECT 0.7950 1.5260 1.6570 1.5760 ;
      RECT 0.2790 0.6180 0.7250 0.6680 ;
      RECT 0.2790 0.6680 0.3290 0.9140 ;
      RECT 0.2790 0.4220 0.3290 0.6180 ;
      RECT 0.7350 0.5180 0.8610 0.5680 ;
      RECT 0.8110 0.5680 0.8610 0.7180 ;
      RECT 0.7350 0.7180 0.8610 0.7680 ;
      RECT 0.7350 0.3940 0.7850 0.5180 ;
      RECT 0.7350 0.7680 0.7850 0.9140 ;
      RECT 1.6470 0.7510 1.7370 0.8010 ;
      RECT 1.6470 0.8010 1.6970 0.9920 ;
      RECT 1.6870 0.6680 1.7370 0.7510 ;
      RECT 1.6870 0.6180 1.9410 0.6680 ;
      RECT 1.6870 0.5680 1.7370 0.6180 ;
      RECT 1.6310 0.5180 1.7370 0.5680 ;
      RECT 2.5620 1.4280 2.7010 1.4780 ;
      RECT 2.5620 1.2700 2.6120 1.4280 ;
      RECT 2.0870 1.2200 2.6120 1.2700 ;
      RECT 1.3430 0.4680 1.3930 0.6180 ;
      RECT 1.3430 0.2820 1.3930 0.4180 ;
      RECT 1.3430 0.6680 1.3930 1.2540 ;
      RECT 1.3430 0.6180 1.6370 0.6680 ;
      RECT 2.1030 0.4680 2.1530 0.7280 ;
      RECT 1.3430 0.4180 2.1530 0.4680 ;
      RECT 2.2380 0.7780 2.2880 1.2200 ;
      RECT 2.1030 0.7280 2.2880 0.7780 ;
      RECT 1.1910 0.2820 1.2410 0.5180 ;
      RECT 1.0390 0.1960 1.0890 0.5180 ;
      RECT 1.1910 0.5680 1.2410 1.2040 ;
      RECT 1.0390 1.2040 1.2410 1.2540 ;
      RECT 1.0390 0.7500 1.0890 1.2040 ;
      RECT 1.0390 0.5180 1.2410 0.5680 ;
      RECT 0.6430 0.0960 1.7890 0.1460 ;
      RECT 1.7070 1.5310 2.0930 1.5810 ;
      RECT 2.0110 0.0960 3.1570 0.1460 ;
    LAYER PO ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 1.2770 0.0680 1.3070 0.6420 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 1.2770 0.9900 1.3070 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 4.3170 0.0680 4.3470 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 2.0370 0.0680 2.0670 0.9060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 2.0370 1.0820 2.0670 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 3.7090 0.0680 3.7390 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
  END
END CGLPPSX4_LVT

MACRO CGLPPSX8_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.016 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.3830 0.1480 4.4330 0.5040 ;
        RECT 3.4710 0.5040 4.8190 0.5530 ;
        RECT 4.6870 0.1480 4.7370 0.5040 ;
        RECT 4.0790 0.1480 4.1290 0.5040 ;
        RECT 3.7750 0.1480 3.8250 0.5040 ;
        RECT 3.4710 0.1480 3.5210 0.5040 ;
        RECT 3.4710 0.5530 4.9190 0.5540 ;
        RECT 4.7690 0.5540 4.9190 0.6630 ;
        RECT 4.7690 0.6630 4.8190 0.8040 ;
        RECT 3.4710 0.8040 4.8190 0.8540 ;
        RECT 4.3830 0.8540 4.4330 1.5460 ;
        RECT 4.6870 0.8540 4.7370 1.5460 ;
        RECT 4.0790 0.8540 4.1290 1.5460 ;
        RECT 3.7750 0.8540 3.8250 1.5460 ;
        RECT 3.4710 0.8540 3.5210 1.5460 ;
    END
    ANTENNADIFFAREA 0.6952 ;
  END GCLK

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 0.8570 0.9670 0.9670 ;
        RECT 0.9170 0.6680 0.9670 0.8570 ;
        RECT 0.9170 0.6180 1.0290 0.6680 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END EN

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2250 0.6180 2.3970 0.6680 ;
        RECT 2.2250 0.5530 2.3350 0.6180 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END SE

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 5.0160 1.7020 ;
        RECT 3.9270 0.9040 3.9770 1.6420 ;
        RECT 3.6230 0.9040 3.6730 1.6420 ;
        RECT 4.2310 0.9040 4.2810 1.6420 ;
        RECT 4.5350 0.9040 4.5850 1.6420 ;
        RECT 0.5830 1.3540 0.6330 1.6420 ;
        RECT 3.1670 1.3660 3.2170 1.6420 ;
        RECT 2.2710 1.3850 2.3210 1.6420 ;
        RECT 0.4310 1.3040 1.5450 1.3540 ;
        RECT 2.6950 1.3160 3.2170 1.3660 ;
        RECT 1.7990 1.3350 2.3210 1.3850 ;
        RECT 0.4310 1.0880 0.4810 1.3040 ;
        RECT 1.4950 0.7500 1.5450 1.3040 ;
        RECT 0.8870 1.0370 0.9370 1.3040 ;
        RECT 0.5830 1.1010 0.6330 1.3040 ;
        RECT 3.1670 1.2660 3.2170 1.3160 ;
        RECT 1.7990 1.1420 1.8490 1.3350 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 5.0160 0.0300 ;
        RECT 3.6230 0.0300 3.6730 0.4540 ;
        RECT 3.9270 0.0300 3.9770 0.4540 ;
        RECT 4.2310 0.0300 4.2810 0.4540 ;
        RECT 4.5350 0.0300 4.5850 0.4540 ;
        RECT 0.4310 0.0300 0.4810 0.1960 ;
        RECT 1.8390 0.0300 1.8890 0.3180 ;
        RECT 0.4310 0.1960 0.9370 0.2460 ;
        RECT 1.4790 0.3180 2.3050 0.3680 ;
        RECT 0.4310 0.2460 0.4810 0.4500 ;
        RECT 0.8870 0.2460 0.9370 0.4500 ;
        RECT 0.5830 0.2460 0.6330 0.4500 ;
        RECT 2.2550 0.3680 2.3050 0.4830 ;
        RECT 2.2550 0.2460 2.3050 0.3180 ;
        RECT 2.2550 0.1960 3.0650 0.2460 ;
        RECT 2.5590 0.2460 2.6090 0.4680 ;
        RECT 3.0150 0.2460 3.0650 0.5820 ;
    END
  END VSS

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 1.4240 0.4210 1.5760 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 5.1310 1.7880 ;
    LAYER M1 ;
      RECT 2.8630 0.7860 3.3090 0.8360 ;
      RECT 2.9030 0.5680 2.9530 0.7860 ;
      RECT 2.8630 0.8360 2.9130 1.1030 ;
      RECT 2.8630 0.5180 2.9530 0.5680 ;
      RECT 2.5420 1.1030 2.9130 1.1530 ;
      RECT 2.8630 0.2960 2.9130 0.5180 ;
      RECT 2.8630 1.1530 2.9130 1.2660 ;
      RECT 2.0110 0.0960 3.1570 0.1460 ;
      RECT 1.0390 1.2040 1.2410 1.2540 ;
      RECT 1.0390 0.7500 1.0890 1.2040 ;
      RECT 1.1910 0.5680 1.2410 1.2040 ;
      RECT 1.0390 0.1960 1.0890 0.5180 ;
      RECT 1.1910 0.2820 1.2410 0.5180 ;
      RECT 1.0390 0.5180 1.2410 0.5680 ;
      RECT 1.6310 0.5180 1.7370 0.5680 ;
      RECT 1.6870 0.5680 1.7370 0.6180 ;
      RECT 1.6870 0.6180 1.9410 0.6680 ;
      RECT 1.6870 0.6680 1.7370 0.7510 ;
      RECT 1.6470 0.7510 1.7370 0.8010 ;
      RECT 1.6470 0.8010 1.6970 0.9920 ;
      RECT 3.3190 0.6040 4.6770 0.6540 ;
      RECT 3.3590 0.6540 3.4090 0.8860 ;
      RECT 3.3190 0.2820 3.3690 0.6040 ;
      RECT 3.3190 0.8860 3.4090 0.9360 ;
      RECT 3.3190 0.9360 3.3690 1.1660 ;
      RECT 3.3190 1.2160 3.3690 1.3580 ;
      RECT 2.9980 1.1660 3.3690 1.2160 ;
      RECT 2.4940 0.6180 2.8530 0.6680 ;
      RECT 2.4940 0.6680 2.5440 0.7200 ;
      RECT 2.4940 0.5680 2.5440 0.6180 ;
      RECT 2.4070 0.7200 2.5440 0.7700 ;
      RECT 2.4070 0.5180 2.5440 0.5680 ;
      RECT 2.4070 0.7700 2.4570 1.1620 ;
      RECT 2.4070 0.3940 2.4570 0.5180 ;
      RECT 1.9760 0.8780 2.0260 1.0420 ;
      RECT 1.9760 0.8280 2.0930 0.8780 ;
      RECT 1.6070 1.0420 2.0260 1.0920 ;
      RECT 1.6070 1.0920 1.6570 1.5260 ;
      RECT 0.7950 1.5260 1.6570 1.5760 ;
      RECT 0.2790 0.6180 0.7250 0.6680 ;
      RECT 0.2790 0.6680 0.3290 0.9140 ;
      RECT 0.2790 0.4220 0.3290 0.6180 ;
      RECT 0.7350 0.5180 0.8610 0.5680 ;
      RECT 0.8110 0.5680 0.8610 0.7180 ;
      RECT 0.7350 0.7180 0.8610 0.7680 ;
      RECT 0.7350 0.3940 0.7850 0.5180 ;
      RECT 0.7350 0.7680 0.7850 0.9140 ;
      RECT 2.5620 1.4280 2.7010 1.4780 ;
      RECT 2.5620 1.2700 2.6120 1.4280 ;
      RECT 2.0870 1.2200 2.6120 1.2700 ;
      RECT 1.3430 0.4680 1.3930 0.6180 ;
      RECT 1.3430 0.2820 1.3930 0.4180 ;
      RECT 1.3430 0.6680 1.3930 1.2540 ;
      RECT 1.3430 0.6180 1.6370 0.6680 ;
      RECT 2.1030 0.4680 2.1530 0.7280 ;
      RECT 1.3430 0.4180 2.1530 0.4680 ;
      RECT 2.2380 0.7780 2.2880 1.2200 ;
      RECT 2.1030 0.7280 2.2880 0.7780 ;
      RECT 0.6430 0.0960 1.7890 0.1460 ;
      RECT 1.7070 1.5310 2.0930 1.5810 ;
    LAYER PO ;
      RECT 2.3410 0.0680 2.3710 1.6060 ;
      RECT 0.0610 0.0680 0.0910 1.6060 ;
      RECT 0.2130 0.0680 0.2430 1.6060 ;
      RECT 2.0370 1.0820 2.0670 1.6060 ;
      RECT 0.8210 0.0680 0.8510 1.6060 ;
      RECT 3.8610 0.0680 3.8910 1.6060 ;
      RECT 2.7970 0.0680 2.8270 1.6060 ;
      RECT 2.1890 0.0680 2.2190 1.6060 ;
      RECT 0.3650 0.0680 0.3950 1.6060 ;
      RECT 2.6450 0.0680 2.6750 1.6060 ;
      RECT 1.8850 0.0680 1.9150 1.6060 ;
      RECT 0.5170 0.0680 0.5470 1.6060 ;
      RECT 2.9490 0.0680 2.9790 1.6060 ;
      RECT 3.7090 0.0680 3.7390 1.6060 ;
      RECT 1.1250 0.0680 1.1550 1.6060 ;
      RECT 0.6690 0.0680 0.6990 1.6060 ;
      RECT 3.5570 0.0680 3.5870 1.6060 ;
      RECT 1.5810 0.0680 1.6110 1.6060 ;
      RECT 3.4050 0.0680 3.4350 1.6060 ;
      RECT 1.2770 0.0680 1.3070 0.6420 ;
      RECT 1.2770 0.9900 1.3070 1.6060 ;
      RECT 2.4930 0.0680 2.5230 1.6060 ;
      RECT 1.7330 0.0680 1.7630 1.6060 ;
      RECT 1.4290 0.0680 1.4590 1.6060 ;
      RECT 2.0370 0.0680 2.0670 0.9060 ;
      RECT 4.0130 0.0680 4.0430 1.6060 ;
      RECT 3.1010 0.0680 3.1310 1.6060 ;
      RECT 4.3170 0.0680 4.3470 1.6060 ;
      RECT 0.9730 0.0680 1.0030 1.6060 ;
      RECT 4.4690 0.0680 4.4990 1.6060 ;
      RECT 4.1650 0.0680 4.1950 1.6060 ;
      RECT 4.7730 0.0680 4.8030 1.6060 ;
      RECT 4.6210 0.0680 4.6510 1.6060 ;
      RECT 4.9250 0.0680 4.9550 1.6060 ;
      RECT 3.2530 0.0680 3.2830 1.6060 ;
  END
END CGLPPSX8_LVT

MACRO AOI21X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.976 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 0.0970 0.8770 0.2070 ;
    END
    ANTENNAGATEAREA 0.0213 ;
  END A3

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.9760 1.7020 ;
        RECT 1.0390 1.0210 1.0890 1.6420 ;
        RECT 0.2790 1.1200 0.3290 1.6420 ;
        RECT 0.5830 1.2120 0.6330 1.6420 ;
        RECT 1.4950 1.2780 1.5450 1.6420 ;
    END
  END VDD

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4910 0.8570 0.6630 0.9670 ;
    END
    ANTENNAGATEAREA 0.0243 ;
  END A1

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.9760 0.0300 ;
        RECT 1.0390 0.0300 1.0890 0.5620 ;
        RECT 1.4950 0.0300 1.5450 0.3970 ;
        RECT 0.2790 0.0300 0.3290 0.2950 ;
        RECT 0.2790 0.2950 0.7850 0.3450 ;
        RECT 0.7350 0.3450 0.7850 0.5690 ;
        RECT 0.2790 0.3450 0.3290 0.5690 ;
    END
  END VSS

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7050 0.4210 0.8150 ;
    END
    ANTENNAGATEAREA 0.0243 ;
  END A2

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6170 1.0090 1.7270 1.1190 ;
        RECT 1.6480 1.1190 1.6980 1.4700 ;
        RECT 1.6480 0.7500 1.6980 1.0090 ;
        RECT 1.6480 0.7000 1.7360 0.7500 ;
        RECT 1.6860 0.5180 1.7360 0.7000 ;
        RECT 1.3190 0.4680 1.7360 0.5180 ;
        RECT 1.3190 0.5180 1.3690 0.7440 ;
        RECT 1.6480 0.1600 1.6980 0.4680 ;
        RECT 1.3430 0.1600 1.3930 0.4680 ;
        RECT 1.3190 0.7440 1.3930 0.7940 ;
        RECT 1.3430 0.7940 1.3930 1.1020 ;
    END
    ANTENNADIFFAREA 0.2484 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 2.0910 1.7870 ;
    LAYER M1 ;
      RECT 1.4190 0.5680 1.6210 0.6500 ;
      RECT 1.1910 1.2020 1.2410 1.5630 ;
      RECT 1.1910 1.0900 1.2410 1.1520 ;
      RECT 1.1910 0.3880 1.2410 0.6060 ;
      RECT 1.1910 1.0400 1.2690 1.0900 ;
      RECT 1.1910 0.6060 1.2690 0.6560 ;
      RECT 1.2190 0.6560 1.2690 1.0400 ;
      RECT 1.4950 0.6500 1.5450 1.1520 ;
      RECT 1.1910 1.1520 1.5450 1.2020 ;
      RECT 1.1170 0.7120 1.1670 0.7760 ;
      RECT 0.8870 0.7760 1.1670 0.8260 ;
      RECT 0.5830 0.3950 0.6330 0.6510 ;
      RECT 0.8870 0.8260 0.9370 1.5750 ;
      RECT 0.8870 0.7010 0.9370 0.7760 ;
      RECT 0.5830 0.6510 0.9370 0.7010 ;
      RECT 0.8870 0.3950 0.9370 0.6510 ;
      RECT 0.7350 1.1270 0.7850 1.5700 ;
      RECT 0.4310 1.0770 0.7850 1.1270 ;
      RECT 0.4310 1.1270 0.4810 1.5750 ;
    LAYER PO ;
      RECT 1.7330 0.0560 1.7630 1.5970 ;
      RECT 0.9730 0.0640 1.0030 1.6130 ;
      RECT 1.1250 0.0590 1.1550 1.6130 ;
      RECT 1.2770 0.0590 1.3070 1.6130 ;
      RECT 0.2130 0.0640 0.2430 1.6130 ;
      RECT 1.4290 0.0640 1.4590 1.6040 ;
      RECT 1.5810 0.0520 1.6110 1.6040 ;
      RECT 0.5170 0.0710 0.5470 1.6200 ;
      RECT 0.0610 0.0640 0.0910 1.6130 ;
      RECT 1.8850 0.0560 1.9150 1.5970 ;
      RECT 0.3650 0.0660 0.3950 1.6200 ;
      RECT 0.6690 0.0710 0.6990 1.6200 ;
      RECT 0.8210 0.0660 0.8510 1.6200 ;
  END
END AOI21X2_LVT

MACRO AOI221X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.128 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7690 1.1610 1.8790 1.2710 ;
        RECT 1.7990 1.2710 1.8490 1.4720 ;
        RECT 1.7990 0.8530 1.8490 1.1610 ;
        RECT 1.7990 0.8520 1.8890 0.8530 ;
        RECT 1.7990 0.8030 1.8990 0.8520 ;
        RECT 1.8490 0.4900 1.8990 0.8030 ;
        RECT 1.7990 0.4260 1.8990 0.4900 ;
        RECT 1.7990 0.1140 1.8490 0.4260 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 0.0970 0.8630 0.2070 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END A3

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.1280 0.0300 ;
        RECT 1.3430 0.0300 1.3930 0.4890 ;
        RECT 1.6470 0.0300 1.6970 0.5110 ;
        RECT 0.5830 0.0300 0.6330 0.4190 ;
        RECT 1.0400 0.0300 1.0900 0.3340 ;
    END
  END VSS

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 0.5530 0.5550 0.6630 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END A2

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.1280 1.7020 ;
        RECT 1.3430 1.1670 1.3930 1.6420 ;
        RECT 0.4310 1.3730 0.4810 1.6420 ;
        RECT 1.6470 1.2060 1.6970 1.6420 ;
    END
  END VDD

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.0090 0.6630 1.1190 ;
        RECT 0.6130 0.9000 0.6630 1.0090 ;
        RECT 0.6130 0.8500 0.7250 0.9000 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END A4

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.8320 0.4040 0.9420 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END A1

  PIN A5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0070 0.7730 1.1810 0.8230 ;
        RECT 1.0090 0.7050 1.1190 0.7730 ;
    END
    ANTENNAGATEAREA 0.0201 ;
  END A5
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 2.2430 1.7870 ;
    LAYER M1 ;
      RECT 1.4190 0.7740 1.4690 0.9070 ;
      RECT 0.8870 0.9070 1.4690 0.9450 ;
      RECT 1.2330 0.9450 1.4690 0.9570 ;
      RECT 0.8870 0.8950 1.2830 0.9070 ;
      RECT 1.2330 0.9570 1.2830 1.0170 ;
      RECT 1.2330 0.7230 1.2830 0.8950 ;
      RECT 1.1910 1.0170 1.2830 1.0810 ;
      RECT 1.1910 1.0810 1.2410 1.5570 ;
      RECT 1.1910 0.6730 1.2820 0.6740 ;
      RECT 1.1910 0.2530 1.2410 0.6730 ;
      RECT 1.1910 0.6740 1.2830 0.7230 ;
      RECT 0.8870 0.7810 0.9370 0.8950 ;
      RECT 0.2790 0.7310 0.9370 0.7810 ;
      RECT 0.8870 0.2620 0.9370 0.7310 ;
      RECT 0.2790 0.2410 0.3290 0.7310 ;
      RECT 1.4950 0.6230 1.7890 0.6730 ;
      RECT 1.6150 0.6730 1.6650 1.0020 ;
      RECT 1.4950 1.0020 1.6650 1.0520 ;
      RECT 1.4950 0.3150 1.5450 0.6230 ;
      RECT 1.4950 1.0520 1.5450 1.5490 ;
      RECT 0.7350 1.0070 1.0890 1.0570 ;
      RECT 1.0390 1.0570 1.0890 1.5570 ;
      RECT 0.7350 1.0570 0.7850 1.2230 ;
      RECT 0.5830 1.3230 0.6330 1.5570 ;
      RECT 0.8870 1.3230 0.9370 1.5570 ;
      RECT 0.2790 1.2730 0.9370 1.3230 ;
      RECT 0.2790 1.3230 0.3290 1.5570 ;
    LAYER PO ;
      RECT 1.8850 0.0630 1.9150 1.6040 ;
      RECT 1.5810 0.0630 1.6110 1.6040 ;
      RECT 1.2770 0.0750 1.3070 1.6210 ;
      RECT 1.7330 0.0640 1.7630 1.6040 ;
      RECT 1.4290 0.0590 1.4590 1.6210 ;
      RECT 2.0370 0.0630 2.0670 1.6040 ;
      RECT 0.6690 0.0720 0.6990 1.6210 ;
      RECT 0.5170 0.0720 0.5470 1.6210 ;
      RECT 0.3650 0.0670 0.3950 1.6210 ;
      RECT 0.0610 0.0720 0.0910 1.6210 ;
      RECT 0.9730 0.0760 1.0030 1.6210 ;
      RECT 0.8210 0.0720 0.8510 1.6210 ;
      RECT 0.2130 0.0720 0.2430 1.6210 ;
      RECT 1.1250 0.0760 1.1550 1.6210 ;
  END
END AOI221X1_LVT

MACRO AOI221X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.28 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9210 1.0090 2.0310 1.1190 ;
        RECT 1.9520 1.1190 2.0020 1.4700 ;
        RECT 1.9520 0.7500 2.0020 1.0090 ;
        RECT 1.9520 0.7000 2.0400 0.7500 ;
        RECT 1.9900 0.5180 2.0400 0.7000 ;
        RECT 1.6230 0.4680 2.0400 0.5180 ;
        RECT 1.6230 0.5180 1.6730 0.7440 ;
        RECT 1.9520 0.1600 2.0020 0.4680 ;
        RECT 1.6470 0.1600 1.6970 0.4680 ;
        RECT 1.6230 0.7440 1.6970 0.7940 ;
        RECT 1.6470 0.7940 1.6970 1.1020 ;
    END
    ANTENNADIFFAREA 0.2484 ;
  END Y

  PIN A5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0070 0.7730 1.1810 0.8230 ;
        RECT 1.0090 0.8230 1.1190 0.8240 ;
        RECT 1.0090 0.7050 1.1190 0.7730 ;
    END
    ANTENNAGATEAREA 0.0228 ;
  END A5

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.8500 0.4300 0.9670 ;
    END
    ANTENNAGATEAREA 0.0252 ;
  END A1

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.0090 0.6630 1.1190 ;
        RECT 0.6130 0.9110 0.6630 1.0090 ;
        RECT 0.6130 0.8610 0.7250 0.9110 ;
    END
    ANTENNAGATEAREA 0.0252 ;
  END A4

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.2800 1.7020 ;
        RECT 1.7990 1.2880 1.8490 1.6420 ;
        RECT 1.3430 1.1120 1.3930 1.6420 ;
        RECT 0.4310 1.3870 0.4810 1.6420 ;
    END
  END VDD

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 0.5530 0.5560 0.6630 ;
    END
    ANTENNAGATEAREA 0.0252 ;
  END A2

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.2800 0.0300 ;
        RECT 1.3430 0.0300 1.3930 0.5130 ;
        RECT 1.7990 0.0300 1.8490 0.3800 ;
        RECT 1.0400 0.0300 1.0900 0.4140 ;
        RECT 0.5830 0.0300 0.6330 0.4370 ;
    END
  END VSS

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 0.0970 0.8630 0.2070 ;
    END
    ANTENNAGATEAREA 0.0252 ;
  END A3
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 2.3950 1.7870 ;
    LAYER M1 ;
      RECT 1.7230 0.5680 1.9250 0.6500 ;
      RECT 1.7990 0.6500 1.8490 1.1700 ;
      RECT 1.4950 1.1700 1.8490 1.2200 ;
      RECT 1.4950 1.2200 1.5450 1.5630 ;
      RECT 1.4950 1.1050 1.5450 1.1700 ;
      RECT 1.4950 0.1550 1.5450 0.6060 ;
      RECT 1.4950 1.0550 1.5730 1.1050 ;
      RECT 1.4950 0.6060 1.5730 0.6560 ;
      RECT 1.5230 0.6560 1.5730 1.0550 ;
      RECT 1.4200 0.8480 1.4700 0.9110 ;
      RECT 0.8870 0.9110 1.4700 0.9580 ;
      RECT 1.1900 0.9580 1.4700 0.9610 ;
      RECT 0.8870 0.7630 0.9370 0.9080 ;
      RECT 0.8870 0.5150 0.9370 0.7130 ;
      RECT 0.8870 0.2610 0.9370 0.4650 ;
      RECT 0.2790 0.7130 0.9370 0.7630 ;
      RECT 0.8870 0.9080 1.2400 0.9110 ;
      RECT 1.1900 0.9610 1.2400 1.4840 ;
      RECT 0.8870 0.5140 1.2260 0.5150 ;
      RECT 0.8870 0.4650 1.2410 0.5140 ;
      RECT 1.1910 0.2400 1.2410 0.4650 ;
      RECT 0.2790 0.2250 0.3290 0.7130 ;
      RECT 1.0390 1.0710 1.0890 1.5700 ;
      RECT 0.7350 1.0250 1.0890 1.0710 ;
      RECT 0.7350 1.0710 0.7850 1.2370 ;
      RECT 0.7550 1.0210 1.0890 1.0250 ;
      RECT 0.8870 1.3370 0.9370 1.5720 ;
      RECT 0.5830 1.3370 0.6330 1.5720 ;
      RECT 0.2790 1.2870 0.9370 1.3370 ;
      RECT 0.2790 1.3370 0.3290 1.5720 ;
    LAYER PO ;
      RECT 2.0370 0.0560 2.0670 1.6190 ;
      RECT 1.7330 0.0640 1.7630 1.6200 ;
      RECT 2.1890 0.0560 2.2190 1.5970 ;
      RECT 1.5810 0.0760 1.6110 1.6210 ;
      RECT 1.2770 0.0760 1.3070 1.6210 ;
      RECT 1.8850 0.0520 1.9150 1.6180 ;
      RECT 1.4290 0.0590 1.4590 1.6130 ;
      RECT 1.1250 0.0770 1.1550 1.6210 ;
      RECT 0.2130 0.0720 0.2430 1.6210 ;
      RECT 0.8210 0.0720 0.8510 1.6210 ;
      RECT 0.9730 0.0760 1.0030 1.6210 ;
      RECT 0.0610 0.0720 0.0910 1.6210 ;
      RECT 0.3650 0.0670 0.3950 1.6210 ;
      RECT 0.5170 0.0720 0.5470 1.6210 ;
      RECT 0.6690 0.0720 0.6990 1.6210 ;
  END
END AOI221X2_LVT

MACRO AOI222X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.28 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9210 1.1610 2.0310 1.2710 ;
        RECT 1.9510 1.2710 2.0010 1.4720 ;
        RECT 1.9510 0.8530 2.0010 1.1610 ;
        RECT 1.9510 0.8520 2.0410 0.8530 ;
        RECT 1.9510 0.8030 2.0510 0.8520 ;
        RECT 2.0010 0.5540 2.0510 0.8030 ;
        RECT 1.9510 0.5040 2.0510 0.5540 ;
        RECT 1.9510 0.1950 2.0010 0.5040 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN A5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0090 0.7690 1.1810 0.8190 ;
        RECT 1.0090 0.6910 1.1190 0.7690 ;
    END
    ANTENNAGATEAREA 0.0228 ;
  END A5

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.8430 0.4040 0.9670 ;
    END
    ANTENNAGATEAREA 0.0228 ;
  END A1

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.0090 0.6630 1.1190 ;
        RECT 0.6130 0.9030 0.6630 1.0090 ;
        RECT 0.6130 0.8530 0.7250 0.9030 ;
    END
    ANTENNAGATEAREA 0.0228 ;
  END A4

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.2800 1.7020 ;
        RECT 1.4950 1.1880 1.5450 1.6420 ;
        RECT 0.4310 1.3730 0.4810 1.6420 ;
        RECT 1.7980 0.7360 1.8480 1.6420 ;
    END
  END VDD

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 0.5530 0.5580 0.6630 ;
    END
    ANTENNAGATEAREA 0.0228 ;
  END A2

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.2800 0.0300 ;
        RECT 1.4950 0.0300 1.5450 0.4860 ;
        RECT 1.7990 0.0300 1.8490 0.5540 ;
        RECT 1.3430 0.0300 1.3930 0.4370 ;
        RECT 0.5830 0.0300 0.6330 0.4650 ;
    END
  END VSS

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 0.0970 0.8630 0.2070 ;
    END
    ANTENNAGATEAREA 0.0228 ;
  END A3

  PIN A6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1590 0.4010 1.2720 0.5110 ;
        RECT 1.1590 0.5110 1.2090 0.5830 ;
        RECT 1.1590 0.5830 1.3330 0.6330 ;
    END
    ANTENNAGATEAREA 0.0228 ;
  END A6
  OBS
    LAYER NWELL ;
      RECT -0.1160 0.6790 2.3960 1.7880 ;
    LAYER M1 ;
      RECT 1.6470 0.6230 1.9410 0.6730 ;
      RECT 1.6470 0.2740 1.6970 0.6230 ;
      RECT 1.6870 0.6730 1.7370 1.0410 ;
      RECT 1.6470 1.0410 1.7370 1.0910 ;
      RECT 1.6470 1.0910 1.6970 1.5630 ;
      RECT 0.8870 0.9080 1.6370 0.9580 ;
      RECT 1.1900 0.9580 1.2400 1.4700 ;
      RECT 1.1900 0.8950 1.2400 0.9080 ;
      RECT 0.2790 0.7750 0.3290 0.7860 ;
      RECT 0.2790 0.2750 0.3290 0.7250 ;
      RECT 0.8870 0.2900 1.0880 0.3400 ;
      RECT 1.0380 0.3400 1.0880 0.4710 ;
      RECT 0.8870 0.7750 0.9370 0.9080 ;
      RECT 0.2790 0.7250 0.9370 0.7750 ;
      RECT 0.8870 0.3400 0.9370 0.7250 ;
      RECT 1.0390 1.5200 1.3920 1.5700 ;
      RECT 1.3420 1.1020 1.3920 1.5200 ;
      RECT 1.0390 1.0990 1.0890 1.5200 ;
      RECT 0.7350 1.0490 1.0890 1.0990 ;
      RECT 0.7350 1.0990 0.7850 1.2230 ;
      RECT 0.8870 1.3230 0.9370 1.5580 ;
      RECT 0.5830 1.3230 0.6330 1.5580 ;
      RECT 0.2790 1.2730 0.9370 1.3230 ;
      RECT 0.2790 1.3230 0.3290 1.5580 ;
    LAYER PO ;
      RECT 2.0370 0.0630 2.0670 1.6040 ;
      RECT 1.7330 0.0630 1.7630 1.6040 ;
      RECT 1.4290 0.0750 1.4590 1.6160 ;
      RECT 1.5810 0.0590 1.6110 1.6130 ;
      RECT 2.1890 0.0630 2.2190 1.6040 ;
      RECT 1.8850 0.0640 1.9150 1.6040 ;
      RECT 1.1250 0.0760 1.1550 1.6210 ;
      RECT 0.2130 0.0720 0.2430 1.6210 ;
      RECT 0.8210 0.0720 0.8510 1.6210 ;
      RECT 0.9730 0.0760 1.0030 1.6210 ;
      RECT 0.0610 0.0720 0.0910 1.6210 ;
      RECT 0.3650 0.0670 0.3950 1.6210 ;
      RECT 0.5170 0.0720 0.5470 1.6210 ;
      RECT 0.6690 0.0720 0.6990 1.6210 ;
      RECT 1.2770 0.0760 1.3070 1.6210 ;
  END
END AOI222X1_LVT

MACRO AOI222X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.432 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0730 1.0090 2.1830 1.1190 ;
        RECT 2.1040 1.1190 2.1540 1.4700 ;
        RECT 2.1040 0.7500 2.1540 1.0090 ;
        RECT 2.1040 0.7000 2.1920 0.7500 ;
        RECT 2.1420 0.5190 2.1920 0.7000 ;
        RECT 1.7750 0.4690 2.1920 0.5190 ;
        RECT 1.7750 0.4680 1.8490 0.4690 ;
        RECT 1.7750 0.5190 1.8250 0.7440 ;
        RECT 2.1030 0.4680 2.1920 0.4690 ;
        RECT 1.7990 0.1600 1.8490 0.4680 ;
        RECT 1.7750 0.7440 1.8490 0.7940 ;
        RECT 2.1030 0.1600 2.1530 0.4680 ;
        RECT 1.7990 0.7940 1.8490 1.1020 ;
    END
    ANTENNADIFFAREA 0.2484 ;
  END Y

  PIN A6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1590 0.4830 1.3330 0.5330 ;
        RECT 1.1590 0.4010 1.2720 0.4830 ;
    END
    ANTENNAGATEAREA 0.0261 ;
  END A6

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 0.0970 0.8630 0.2070 ;
    END
    ANTENNAGATEAREA 0.0261 ;
  END A3

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 0.2490 0.5110 0.3590 ;
        RECT 0.4010 0.3590 0.4510 0.4810 ;
        RECT 0.4010 0.4810 0.5730 0.5310 ;
    END
    ANTENNAGATEAREA 0.0261 ;
  END A2

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 0.9950 0.6630 1.1190 ;
        RECT 0.6130 0.8510 0.6630 0.9950 ;
        RECT 0.6130 0.8010 0.7250 0.8510 ;
    END
    ANTENNAGATEAREA 0.0261 ;
  END A4

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.8430 0.4040 0.9670 ;
        RECT 0.3540 0.7840 0.4040 0.8430 ;
    END
    ANTENNAGATEAREA 0.0261 ;
  END A1

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.4320 0.0300 ;
        RECT 1.9510 0.0300 2.0010 0.3190 ;
        RECT 1.4950 0.0300 1.5450 0.4680 ;
        RECT 0.5830 0.0300 0.6330 0.4000 ;
        RECT 1.3430 0.0300 1.3930 0.4010 ;
    END
  END VSS

  PIN A5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0090 0.7050 1.1190 0.7660 ;
        RECT 1.0090 0.7660 1.1810 0.8160 ;
    END
    ANTENNAGATEAREA 0.0261 ;
  END A5

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.4320 1.7020 ;
        RECT 1.4950 1.1790 1.5450 1.6420 ;
        RECT 1.9510 1.3700 2.0010 1.6420 ;
        RECT 0.4310 1.3730 0.4810 1.6420 ;
    END
  END VDD
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 2.5470 1.7870 ;
    LAYER M1 ;
      RECT 1.8750 0.5730 2.0770 0.6500 ;
      RECT 1.8750 0.6500 2.0540 0.6550 ;
      RECT 1.9510 0.6550 2.0010 1.2290 ;
      RECT 1.6470 1.2290 2.0010 1.2790 ;
      RECT 1.6470 1.2790 1.6970 1.5630 ;
      RECT 1.6470 1.1050 1.6970 1.2290 ;
      RECT 1.6470 0.2600 1.6970 0.6060 ;
      RECT 1.6470 1.0550 1.7250 1.1050 ;
      RECT 1.6470 0.6060 1.7250 0.6560 ;
      RECT 1.6750 0.6560 1.7250 1.0550 ;
      RECT 1.3430 1.0100 1.3930 1.5200 ;
      RECT 1.0390 1.5200 1.3930 1.5700 ;
      RECT 1.0390 1.0990 1.0890 1.5200 ;
      RECT 0.7350 1.0490 1.0890 1.0990 ;
      RECT 0.7350 1.0990 0.7850 1.2230 ;
      RECT 0.8870 0.9080 1.6210 0.9580 ;
      RECT 1.5710 0.8460 1.6210 0.9080 ;
      RECT 0.2790 0.2520 0.3290 0.5840 ;
      RECT 1.1900 0.9580 1.2400 1.4700 ;
      RECT 1.1900 0.8940 1.2400 0.9080 ;
      RECT 0.8870 0.2640 1.0890 0.3130 ;
      RECT 0.9040 0.2630 1.0890 0.2640 ;
      RECT 1.0390 0.3130 1.0890 0.4400 ;
      RECT 0.8870 0.6340 0.9370 0.9080 ;
      RECT 0.2790 0.5840 0.9370 0.6340 ;
      RECT 0.8870 0.3130 0.9370 0.5840 ;
      RECT 0.5830 1.3230 0.6330 1.5580 ;
      RECT 0.8870 1.3230 0.9370 1.5570 ;
      RECT 0.2790 1.2730 0.9370 1.3230 ;
      RECT 0.2790 1.3230 0.3290 1.5570 ;
    LAYER PO ;
      RECT 2.1890 0.0560 2.2190 1.5970 ;
      RECT 1.4290 0.0750 1.4590 1.6160 ;
      RECT 1.8850 0.0640 1.9150 1.6040 ;
      RECT 2.3410 0.0560 2.3710 1.5970 ;
      RECT 2.0370 0.0520 2.0670 1.6040 ;
      RECT 1.2770 0.0760 1.3070 1.6210 ;
      RECT 0.6690 0.0720 0.6990 1.6210 ;
      RECT 0.5170 0.0720 0.5470 1.6210 ;
      RECT 0.3650 0.0670 0.3950 1.6210 ;
      RECT 1.7330 0.0590 1.7630 1.6130 ;
      RECT 0.0610 0.0720 0.0910 1.6210 ;
      RECT 0.9730 0.0760 1.0030 1.6210 ;
      RECT 1.5810 0.0590 1.6110 1.6130 ;
      RECT 0.8210 0.0720 0.8510 1.6210 ;
      RECT 0.2130 0.0720 0.2430 1.6210 ;
      RECT 1.1250 0.0760 1.1550 1.6210 ;
  END
END AOI222X2_LVT

MACRO AOI22X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.824 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4650 1.1610 1.5750 1.2710 ;
        RECT 1.4950 1.2710 1.5450 1.4730 ;
        RECT 1.4950 0.8540 1.5450 1.1610 ;
        RECT 1.4950 0.8040 1.5850 0.8540 ;
        RECT 1.5350 0.4930 1.5850 0.8040 ;
        RECT 1.4950 0.4430 1.5850 0.4930 ;
        RECT 1.4950 0.1350 1.5450 0.4430 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7050 0.4040 0.8150 ;
    END
    ANTENNAGATEAREA 0.0234 ;
  END A1

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 0.5530 0.7080 0.6630 ;
    END
    ANTENNAGATEAREA 0.0234 ;
  END A4

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.8240 1.7020 ;
        RECT 0.4310 1.3710 0.4810 1.6420 ;
        RECT 1.0390 1.0510 1.0890 1.6420 ;
        RECT 1.3420 1.1610 1.3920 1.6420 ;
    END
  END VDD

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 0.0970 0.8630 0.2070 ;
    END
    ANTENNAGATEAREA 0.0234 ;
  END A3

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5070 0.9120 0.5570 1.0090 ;
        RECT 0.4010 1.0090 0.5570 1.1190 ;
    END
    ANTENNAGATEAREA 0.0234 ;
  END A2

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.8240 0.0300 ;
        RECT 1.3430 0.0300 1.3930 0.4730 ;
        RECT 0.5830 0.0300 0.6330 0.3770 ;
        RECT 1.0390 0.0300 1.0890 0.5630 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.9390 1.7870 ;
    LAYER M1 ;
      RECT 1.1910 0.6120 1.4850 0.6620 ;
      RECT 1.3460 0.6620 1.3960 1.0030 ;
      RECT 1.1910 1.0030 1.3960 1.0530 ;
      RECT 1.1910 0.6620 1.2410 0.6630 ;
      RECT 1.1910 0.3890 1.2410 0.6120 ;
      RECT 1.1910 1.0530 1.2410 1.5640 ;
      RECT 1.1910 1.0020 1.2410 1.0030 ;
      RECT 0.8870 1.3210 0.9370 1.5550 ;
      RECT 0.5830 1.3210 0.6330 1.5550 ;
      RECT 0.2790 1.2710 0.9370 1.3210 ;
      RECT 0.2790 1.3210 0.3290 1.5550 ;
      RECT 0.7350 0.8460 1.1810 0.8960 ;
      RECT 0.2790 0.2790 0.3290 0.4520 ;
      RECT 0.7350 0.8130 0.8080 0.8460 ;
      RECT 0.7350 0.8960 0.7850 1.2120 ;
      RECT 0.2790 0.4520 0.9370 0.5020 ;
      RECT 0.8870 0.2790 0.9370 0.4520 ;
      RECT 0.7580 0.5020 0.8080 0.8130 ;
    LAYER PO ;
      RECT 1.5810 0.0640 1.6110 1.6050 ;
      RECT 1.4290 0.0650 1.4590 1.6050 ;
      RECT 0.2130 0.0720 0.2430 1.6210 ;
      RECT 0.8210 0.0720 0.8510 1.6210 ;
      RECT 1.7330 0.0640 1.7630 1.6050 ;
      RECT 0.9730 0.0760 1.0030 1.6210 ;
      RECT 1.2770 0.0600 1.3070 1.6140 ;
      RECT 0.0610 0.0720 0.0910 1.6210 ;
      RECT 0.3650 0.0670 0.3950 1.6210 ;
      RECT 0.5170 0.0720 0.5470 1.6210 ;
      RECT 0.6690 0.0720 0.6990 1.6210 ;
      RECT 1.1250 0.0600 1.1550 1.6140 ;
  END
END AOI22X1_LVT

MACRO AOI22X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.976 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 0.0970 0.8630 0.2270 ;
    END
    ANTENNAGATEAREA 0.0225 ;
  END A3

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2480 0.7050 0.4040 0.8150 ;
    END
    ANTENNAGATEAREA 0.0225 ;
  END A1

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.9760 0.0300 ;
        RECT 0.5830 0.0300 0.6330 0.3640 ;
        RECT 1.0390 0.0300 1.0890 0.4500 ;
        RECT 1.4950 0.0300 1.5450 0.3150 ;
    END
  END VSS

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5070 0.7240 0.5570 1.0090 ;
        RECT 0.4010 1.0090 0.5570 1.1190 ;
    END
    ANTENNAGATEAREA 0.0225 ;
  END A2

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.9760 1.7020 ;
        RECT 0.4310 1.3730 0.4810 1.6420 ;
        RECT 1.0390 1.0210 1.0890 1.6420 ;
        RECT 1.4950 1.3700 1.5450 1.6420 ;
    END
  END VDD

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 0.5530 0.7080 0.6630 ;
    END
    ANTENNAGATEAREA 0.0225 ;
  END A4

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6170 1.0090 1.7270 1.1190 ;
        RECT 1.6480 1.1190 1.6980 1.4700 ;
        RECT 1.6480 0.7500 1.6980 1.0090 ;
        RECT 1.6480 0.7000 1.7360 0.7500 ;
        RECT 1.6860 0.5180 1.7360 0.7000 ;
        RECT 1.3190 0.4680 1.7360 0.5180 ;
        RECT 1.3190 0.5180 1.3690 0.7440 ;
        RECT 1.6480 0.1600 1.6980 0.4680 ;
        RECT 1.3430 0.1600 1.3930 0.4680 ;
        RECT 1.3190 0.7440 1.3930 0.7940 ;
        RECT 1.3430 0.7940 1.3930 1.1020 ;
    END
    ANTENNADIFFAREA 0.2484 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 2.0910 1.7870 ;
    LAYER M1 ;
      RECT 1.4190 0.5680 1.6210 0.6500 ;
      RECT 1.1910 1.2790 1.2410 1.5630 ;
      RECT 1.1910 1.1050 1.2410 1.2290 ;
      RECT 1.1910 0.1840 1.2410 0.6060 ;
      RECT 1.1910 1.0550 1.2690 1.1050 ;
      RECT 1.1910 0.6060 1.2690 0.6560 ;
      RECT 1.2190 0.6560 1.2690 1.0550 ;
      RECT 1.4950 0.6500 1.5450 1.2290 ;
      RECT 1.1910 1.2290 1.5450 1.2790 ;
      RECT 1.1160 0.7120 1.1660 0.8130 ;
      RECT 0.7350 0.8130 1.1660 0.8630 ;
      RECT 0.7350 0.8630 0.7850 1.2230 ;
      RECT 0.2790 0.4420 0.9370 0.4920 ;
      RECT 0.8870 0.2840 0.9370 0.4420 ;
      RECT 0.7580 0.4920 0.8080 0.8130 ;
      RECT 0.2790 0.2810 0.3290 0.4420 ;
      RECT 0.5830 1.3230 0.6330 1.5570 ;
      RECT 0.8870 1.3230 0.9370 1.5570 ;
      RECT 0.2790 1.2730 0.9370 1.3230 ;
      RECT 0.2790 1.3230 0.3290 1.5570 ;
    LAYER PO ;
      RECT 1.7330 0.0560 1.7630 1.5970 ;
      RECT 0.6690 0.0770 0.6990 1.6210 ;
      RECT 0.5170 0.0770 0.5470 1.6210 ;
      RECT 0.3650 0.0720 0.3950 1.6210 ;
      RECT 0.0610 0.0720 0.0910 1.6210 ;
      RECT 0.9730 0.0760 1.0030 1.6210 ;
      RECT 0.8210 0.0770 0.8510 1.6210 ;
      RECT 0.2130 0.0720 0.2430 1.6210 ;
      RECT 1.2770 0.0760 1.3070 1.6210 ;
      RECT 1.5810 0.0520 1.6110 1.6040 ;
      RECT 1.8850 0.0560 1.9150 1.5970 ;
      RECT 1.4290 0.0640 1.4590 1.6040 ;
      RECT 1.1250 0.0590 1.1550 1.6130 ;
  END
END AOI22X2_LVT

MACRO AOINVX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.28 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1570 0.6730 1.3330 0.7330 ;
        RECT 1.1610 0.7330 1.2710 0.8150 ;
    END
    ANTENNAGATEAREA 0.0333 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3430 0.7890 1.5380 0.8390 ;
        RECT 1.3430 0.8390 1.3930 1.5640 ;
        RECT 1.4880 0.6630 1.5380 0.7890 ;
        RECT 1.4650 0.6090 1.5750 0.6630 ;
        RECT 1.3430 0.5590 1.5750 0.6090 ;
        RECT 1.3430 0.2990 1.3930 0.5590 ;
        RECT 1.4650 0.5530 1.5750 0.5590 ;
    END
    ANTENNADIFFAREA 0.1132 ;
  END Y

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.8180 1.0090 1.0080 1.1190 ;
        RECT 0.8820 0.9910 0.9420 1.0090 ;
        RECT 0.8820 1.1190 0.9420 1.2830 ;
        RECT 0.8820 1.2830 1.2410 1.3330 ;
        RECT 1.1910 1.3330 1.2410 1.5640 ;
        RECT 1.1910 0.9300 1.2410 1.2830 ;
    END
  END VDDG

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.2800 1.7020 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.2800 0.0300 ;
        RECT 1.1910 0.0300 1.2410 0.6090 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 2.2800 3.3740 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT 0.7990 0.6790 1.5920 2.6650 ;
    LAYER PO ;
      RECT 1.2770 1.7390 1.3070 3.2340 ;
      RECT 0.5170 1.7390 0.5470 3.2340 ;
      RECT 1.4290 1.7390 1.4590 3.2340 ;
      RECT 1.5810 1.7390 1.6110 3.2340 ;
      RECT 0.8210 1.7390 0.8510 3.2340 ;
      RECT 0.2130 1.7390 0.2430 3.2340 ;
      RECT 0.3650 1.7390 0.3950 3.2340 ;
      RECT 0.9730 1.7390 1.0030 3.2340 ;
      RECT 0.6690 1.7390 0.6990 3.2340 ;
      RECT 1.7330 1.7390 1.7630 3.2340 ;
      RECT 1.8850 1.7390 1.9150 3.2340 ;
      RECT 0.6690 0.1120 0.6990 1.6240 ;
      RECT 0.5170 0.1120 0.5470 1.6240 ;
      RECT 0.3650 0.1120 0.3950 1.6240 ;
      RECT 0.2130 0.1120 0.2430 1.6240 ;
      RECT 1.8850 0.1120 1.9150 1.6240 ;
      RECT 1.7330 0.1120 1.7630 1.6240 ;
      RECT 1.5810 0.1120 1.6110 1.6240 ;
      RECT 2.0370 1.7390 2.0670 3.2340 ;
      RECT 2.0370 0.1120 2.0670 1.6240 ;
      RECT 2.1890 1.7390 2.2190 3.2340 ;
      RECT 2.1890 0.1120 2.2190 1.6240 ;
      RECT 0.8210 0.1120 0.8510 1.6240 ;
      RECT 0.0610 1.7390 0.0910 3.2340 ;
      RECT 0.0610 0.1120 0.0910 1.6240 ;
      RECT 0.9730 0.1120 1.0030 1.6240 ;
      RECT 1.1250 0.1120 1.1550 1.6240 ;
      RECT 1.1250 1.7390 1.1550 3.2340 ;
      RECT 1.2770 0.1120 1.3070 1.6240 ;
      RECT 1.4290 0.1120 1.4590 1.6240 ;
  END
END AOINVX1_LVT

MACRO AOINVX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.28 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0050 0.6730 1.3330 0.7330 ;
        RECT 1.0090 0.7330 1.1190 0.8150 ;
    END
    ANTENNAGATEAREA 0.0666 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1910 0.5590 1.5740 0.6090 ;
        RECT 1.1910 0.2990 1.2410 0.5590 ;
        RECT 1.4640 0.6090 1.5740 0.6630 ;
        RECT 1.4640 0.5530 1.5740 0.5590 ;
        RECT 1.4640 0.6630 1.5140 0.7930 ;
        RECT 1.1750 0.7930 1.5140 0.8430 ;
    END
    ANTENNADIFFAREA 0.1354 ;
  END Y

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.6660 1.0090 0.8560 1.1190 ;
        RECT 0.7300 0.9910 0.7900 1.0090 ;
        RECT 0.7300 1.1190 0.7900 1.2430 ;
        RECT 0.7300 1.2430 1.3930 1.2930 ;
        RECT 1.3430 1.2930 1.3930 1.5640 ;
        RECT 1.3430 0.9300 1.3930 1.2430 ;
        RECT 1.0390 1.2930 1.0890 1.5640 ;
        RECT 1.0390 0.9300 1.0890 1.2430 ;
    END
  END VDDG

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.2800 1.7020 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.2800 0.0300 ;
        RECT 1.0390 0.0300 1.0890 0.6090 ;
        RECT 1.3430 0.0300 1.3930 0.5010 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 2.2800 3.3740 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT 0.6280 0.6790 1.6240 2.6650 ;
    LAYER PO ;
      RECT 1.4290 0.2390 1.4590 1.6240 ;
      RECT 1.4290 1.7940 1.4590 3.1790 ;
      RECT 0.6690 1.7940 0.6990 3.1790 ;
      RECT 0.8210 1.7940 0.8510 3.1790 ;
      RECT 0.9730 1.7940 1.0030 3.1790 ;
      RECT 1.5810 1.7940 1.6110 3.1790 ;
      RECT 1.1250 1.7940 1.1550 3.1790 ;
      RECT 1.2770 1.7940 1.3070 3.1790 ;
      RECT 2.0370 1.7940 2.0670 3.1790 ;
      RECT 2.1890 1.7940 2.2190 3.1790 ;
      RECT 1.7330 1.7940 1.7630 3.1790 ;
      RECT 1.8850 1.7940 1.9150 3.1790 ;
      RECT 0.0610 1.7940 0.0910 3.1790 ;
      RECT 0.2130 1.7940 0.2430 3.1790 ;
      RECT 0.3650 1.7940 0.3950 3.1790 ;
      RECT 0.5170 1.7940 0.5470 3.1790 ;
      RECT 0.0610 0.2330 0.0910 1.6180 ;
      RECT 0.2130 0.2330 0.2430 1.6180 ;
      RECT 0.3650 0.2330 0.3950 1.6180 ;
      RECT 0.5170 0.2330 0.5470 1.6180 ;
      RECT 2.0370 0.2390 2.0670 1.6240 ;
      RECT 2.1890 0.2390 2.2190 1.6240 ;
      RECT 1.7330 0.2390 1.7630 1.6240 ;
      RECT 1.8850 0.2390 1.9150 1.6240 ;
      RECT 0.6690 0.2390 0.6990 1.6240 ;
      RECT 0.8210 0.2390 0.8510 1.6240 ;
      RECT 0.9730 0.2390 1.0030 1.6240 ;
      RECT 1.5810 0.2390 1.6110 1.6240 ;
      RECT 1.1250 0.2390 1.1550 1.6240 ;
      RECT 1.2770 0.2390 1.3070 1.6240 ;
  END
END AOINVX2_LVT

MACRO AOINVX4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.584 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0050 0.6730 1.6370 0.7330 ;
        RECT 1.0090 0.7330 1.1190 0.8150 ;
    END
    ANTENNAGATEAREA 0.1332 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1910 0.1890 1.2410 0.5370 ;
        RECT 1.1910 0.5370 1.8750 0.5530 ;
        RECT 1.1910 0.5530 1.8790 0.5870 ;
        RECT 1.4950 0.1890 1.5450 0.5370 ;
        RECT 1.7690 0.5870 1.8790 0.6630 ;
        RECT 1.7690 0.6630 1.8190 0.9250 ;
        RECT 1.1910 0.9250 1.8190 0.9750 ;
        RECT 1.4950 0.9750 1.5450 1.4580 ;
        RECT 1.4950 0.8240 1.5450 0.9250 ;
        RECT 1.1910 0.9750 1.2410 1.4580 ;
        RECT 1.1910 0.8240 1.2410 0.9250 ;
    END
    ANTENNADIFFAREA 0.2708 ;
  END Y

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.6660 1.0090 0.8560 1.1190 ;
        RECT 0.7300 0.9910 0.7900 1.0090 ;
        RECT 0.7300 1.1190 0.7900 1.5080 ;
        RECT 0.7300 1.5080 1.7130 1.5330 ;
        RECT 0.7350 1.5330 1.7130 1.5580 ;
    END
  END VDDG

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.5840 1.7020 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.5840 0.0300 ;
        RECT 1.0390 0.0300 1.0890 0.4530 ;
        RECT 1.3430 0.0300 1.3930 0.4530 ;
        RECT 1.6470 0.0300 1.6970 0.4530 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 2.5840 3.3740 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT 0.6490 0.6790 1.9250 2.6650 ;
    LAYER PO ;
      RECT 1.4290 0.1290 1.4590 1.6240 ;
      RECT 1.5810 0.1290 1.6110 1.6240 ;
      RECT 1.4290 1.7590 1.4590 3.2540 ;
      RECT 1.5810 1.7590 1.6110 3.2540 ;
      RECT 0.6690 1.7590 0.6990 3.2540 ;
      RECT 0.8210 1.7590 0.8510 3.2540 ;
      RECT 1.7330 1.7590 1.7630 3.2540 ;
      RECT 0.9730 1.7590 1.0030 3.2540 ;
      RECT 1.8850 1.7590 1.9150 3.2540 ;
      RECT 1.1250 1.7590 1.1550 3.2540 ;
      RECT 1.2770 1.7590 1.3070 3.2540 ;
      RECT 2.0370 1.7590 2.0670 3.2540 ;
      RECT 2.1890 1.7590 2.2190 3.2540 ;
      RECT 2.3410 1.7590 2.3710 3.2540 ;
      RECT 0.0610 1.7590 0.0910 3.2540 ;
      RECT 0.2130 1.7590 0.2430 3.2540 ;
      RECT 0.3650 1.7590 0.3950 3.2540 ;
      RECT 0.5170 1.7590 0.5470 3.2540 ;
      RECT 0.5170 0.1290 0.5470 1.6240 ;
      RECT 0.3650 0.1290 0.3950 1.6240 ;
      RECT 0.2130 0.1290 0.2430 1.6240 ;
      RECT 0.0610 0.1290 0.0910 1.6240 ;
      RECT 2.3410 0.1290 2.3710 1.6240 ;
      RECT 2.1890 0.1290 2.2190 1.6240 ;
      RECT 0.6690 0.1290 0.6990 1.6240 ;
      RECT 2.0370 0.1290 2.0670 1.6240 ;
      RECT 2.4930 1.7590 2.5230 3.2540 ;
      RECT 0.8210 0.1290 0.8510 1.6240 ;
      RECT 2.4930 0.1290 2.5230 1.6240 ;
      RECT 1.7330 0.1290 1.7630 1.6240 ;
      RECT 0.9730 0.1290 1.0030 1.6240 ;
      RECT 1.8850 0.1290 1.9150 1.6240 ;
      RECT 1.1250 0.1290 1.1550 1.6240 ;
      RECT 1.2770 0.1290 1.3070 1.6240 ;
  END
END AOINVX4_LVT

MACRO BSLEX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.064 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.0640 1.7020 ;
        RECT 0.2790 0.7770 0.3290 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.0640 0.0300 ;
        RECT 0.2240 0.0300 0.2740 0.3590 ;
        RECT 0.2240 0.3590 0.3290 0.4090 ;
        RECT 0.2790 0.4090 0.3290 0.5630 ;
    END
  END VSS

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3240 0.0920 0.7400 0.1420 ;
        RECT 0.3980 0.1420 0.5110 0.2070 ;
    END
    ANTENNAGATEAREA 0.02205 ;
  END EN

  PIN INOUT1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 0.5530 0.6630 0.6630 ;
        RECT 0.5830 0.6630 0.6330 1.4720 ;
        RECT 0.5830 0.1920 0.6330 0.5530 ;
    END
    ANTENNADIFFAREA 0.1111 ;
    ANTENNAGATEAREA 0.1111 ;
  END INOUT1

  PIN INOUT2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 0.7050 0.8150 0.8150 ;
        RECT 0.7350 0.8150 0.7850 1.4720 ;
        RECT 0.7350 0.1920 0.7850 0.7050 ;
    END
    ANTENNADIFFAREA 0.1111 ;
    ANTENNAGATEAREA 0.1111 ;
  END INOUT2
  OBS
    LAYER NWELL ;
      RECT -0.1120 0.6790 1.1760 1.7730 ;
    LAYER M1 ;
      RECT 0.4310 1.5280 0.7400 1.5780 ;
      RECT 0.4310 0.4700 0.4810 1.5780 ;
      RECT 0.4310 0.4200 0.4810 0.4700 ;
    LAYER PO ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.6690 0.7170 0.6990 1.6060 ;
      RECT 0.6690 0.0640 0.6990 0.6150 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
      RECT 0.8210 0.0660 0.8510 1.6060 ;
  END
END BSLEX1_LVT

MACRO BSLEX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.216 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.2160 1.7020 ;
        RECT 0.2790 0.7770 0.3290 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.2160 0.0300 ;
        RECT 0.2240 0.0300 0.2740 0.1920 ;
        RECT 0.2240 0.1920 0.3290 0.2420 ;
        RECT 0.2790 0.2420 0.3290 0.5630 ;
    END
  END VSS

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3240 0.0920 1.1190 0.1420 ;
        RECT 1.0090 0.1420 1.1190 0.2070 ;
    END
    ANTENNAGATEAREA 0.0387 ;
  END EN

  PIN INOUT1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5330 0.5530 0.6630 0.6630 ;
        RECT 0.5830 0.6630 0.6330 1.4220 ;
        RECT 0.5830 0.1920 0.6330 0.5530 ;
        RECT 0.5830 1.4220 0.9370 1.4720 ;
        RECT 0.8870 0.1920 0.9370 1.4220 ;
    END
    ANTENNADIFFAREA 0.2222 ;
    ANTENNAGATEAREA 0.2222 ;
  END INOUT1

  PIN INOUT2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 1.1600 0.8370 1.2710 ;
        RECT 0.7350 1.2710 0.7850 1.2880 ;
        RECT 0.7350 0.1920 0.7850 1.1600 ;
    END
    ANTENNADIFFAREA 0.133 ;
    ANTENNAGATEAREA 0.133 ;
  END INOUT2
  OBS
    LAYER NWELL ;
      RECT -0.1120 0.6790 1.3280 1.7730 ;
    LAYER M1 ;
      RECT 0.4310 1.5280 0.8920 1.5780 ;
      RECT 0.4310 0.4170 0.4810 1.5780 ;
      RECT 0.4310 0.3670 0.4810 0.4170 ;
      RECT 0.4310 0.3590 0.4810 0.4170 ;
    LAYER PO ;
      RECT 0.6690 0.0660 0.6990 0.6150 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 0.8210 0.0660 0.8510 0.6150 ;
      RECT 0.8210 0.7170 0.8510 1.6060 ;
      RECT 1.1250 0.0660 1.1550 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.6690 0.7170 0.6990 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
      RECT 0.9730 0.0660 1.0030 1.6060 ;
  END
END BSLEX2_LVT

MACRO BSLEX4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.52 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.5200 1.7020 ;
        RECT 0.2790 0.7770 0.3290 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.5200 0.0300 ;
        RECT 0.2240 0.0300 0.2740 0.1920 ;
        RECT 0.2240 0.1920 0.3290 0.2420 ;
        RECT 0.2790 0.2420 0.3290 0.5630 ;
    END
  END VSS

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3240 0.0920 1.4210 0.0950 ;
        RECT 0.3240 0.0950 1.4230 0.1420 ;
        RECT 1.3110 0.1420 1.4230 0.2070 ;
    END
    ANTENNAGATEAREA 0.0777 ;
  END EN

  PIN INOUT1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 0.5530 0.6630 0.6630 ;
        RECT 0.5830 0.6630 0.6330 1.4220 ;
        RECT 0.5830 0.1920 0.6330 0.5530 ;
        RECT 0.5830 1.4220 1.2410 1.4720 ;
        RECT 0.8870 0.3250 0.9370 1.4220 ;
        RECT 1.1910 0.1920 1.2410 1.4220 ;
    END
    ANTENNADIFFAREA 0.3552 ;
    ANTENNAGATEAREA 0.3552 ;
  END INOUT1

  PIN INOUT2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 1.1600 0.8350 1.2710 ;
        RECT 0.7350 1.2710 0.7850 1.2880 ;
        RECT 0.7350 0.2420 0.7850 1.1600 ;
        RECT 0.7350 0.1920 1.0890 0.2420 ;
        RECT 1.0390 0.2420 1.0890 1.2880 ;
    END
    ANTENNADIFFAREA 0.266 ;
    ANTENNAGATEAREA 0.266 ;
  END INOUT2
  OBS
    LAYER NWELL ;
      RECT -0.1120 0.6790 1.6320 1.7730 ;
    LAYER M1 ;
      RECT 0.4310 1.5280 1.1960 1.5780 ;
      RECT 0.4310 0.3220 0.4810 1.5780 ;
      RECT 0.4310 0.2720 0.4810 0.3220 ;
    LAYER PO ;
      RECT 1.1250 0.0660 1.1550 0.6150 ;
      RECT 1.1250 0.7170 1.1550 1.6060 ;
      RECT 0.9730 0.0660 1.0030 0.6150 ;
      RECT 0.9730 0.7170 1.0030 1.6060 ;
      RECT 0.6690 0.0660 0.6990 0.6150 ;
      RECT 1.4290 0.0660 1.4590 1.6060 ;
      RECT 0.2130 0.0660 0.2430 1.6060 ;
      RECT 0.8210 0.0660 0.8510 0.6150 ;
      RECT 0.8210 0.7170 0.8510 1.6060 ;
      RECT 1.2770 0.0660 1.3070 1.6060 ;
      RECT 0.0610 0.0660 0.0910 1.6060 ;
      RECT 0.6690 0.7170 0.6990 1.6060 ;
      RECT 0.5170 0.0660 0.5470 1.6060 ;
      RECT 0.3650 0.0660 0.3950 1.6060 ;
  END
END BSLEX4_LVT

MACRO AO221X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.976 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.9760 0.0300 ;
        RECT 1.4950 0.0300 1.5450 0.3940 ;
        RECT 0.5830 0.0300 0.6330 0.3660 ;
        RECT 1.0400 0.0300 1.0900 0.3970 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6170 1.0090 1.7270 1.1190 ;
        RECT 1.6480 1.1190 1.6980 1.4700 ;
        RECT 1.6480 0.7830 1.6980 1.0090 ;
        RECT 1.6480 0.7330 1.7360 0.7830 ;
        RECT 1.6860 0.5530 1.7360 0.7330 ;
        RECT 1.3150 0.5030 1.7360 0.5530 ;
        RECT 1.3150 0.5530 1.3650 0.7440 ;
        RECT 1.6480 0.4820 1.7360 0.5030 ;
        RECT 1.3430 0.1740 1.3930 0.5030 ;
        RECT 1.3150 0.7440 1.3930 0.8060 ;
        RECT 1.6480 0.1740 1.6980 0.4820 ;
        RECT 1.3430 0.8060 1.3930 1.1020 ;
    END
    ANTENNADIFFAREA 0.2484 ;
  END Y

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 0.0970 0.8630 0.2070 ;
    END
    ANTENNAGATEAREA 0.0279 ;
  END A3

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 0.2490 0.5110 0.3590 ;
        RECT 0.4010 0.3590 0.4510 0.4980 ;
        RECT 0.4010 0.4980 0.5730 0.5480 ;
    END
    ANTENNAGATEAREA 0.0279 ;
  END A2

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.9760 1.7020 ;
        RECT 1.4950 1.2700 1.5450 1.6420 ;
        RECT 0.4310 1.3730 0.4810 1.6420 ;
    END
  END VDD

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.0090 0.6630 1.1190 ;
        RECT 0.6060 0.8080 0.6560 1.0090 ;
        RECT 0.6060 0.7580 0.7250 0.8080 ;
    END
    ANTENNAGATEAREA 0.0279 ;
  END A4

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.8570 0.4050 0.9670 ;
        RECT 0.3550 0.7350 0.4050 0.8570 ;
    END
    ANTENNAGATEAREA 0.0279 ;
  END A1

  PIN A5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0090 0.7050 1.1190 0.7590 ;
        RECT 1.0090 0.7590 1.1810 0.8090 ;
        RECT 1.0090 0.8090 1.1190 0.8150 ;
    END
    ANTENNAGATEAREA 0.0246 ;
  END A5
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 2.0910 1.7730 ;
    LAYER M1 ;
      RECT 1.4190 0.6030 1.6210 0.6830 ;
      RECT 1.4190 0.6830 1.5980 0.6850 ;
      RECT 1.4930 0.6850 1.5430 1.1700 ;
      RECT 1.1900 1.1700 1.5430 1.2200 ;
      RECT 1.1900 1.2200 1.2400 1.5570 ;
      RECT 1.1900 0.9670 1.2400 1.1700 ;
      RECT 0.8870 0.9170 1.2400 0.9670 ;
      RECT 0.8870 0.5820 1.2420 0.5980 ;
      RECT 1.1920 0.3090 1.2420 0.5820 ;
      RECT 0.2790 0.5980 1.2420 0.6320 ;
      RECT 0.8870 0.6480 0.9370 0.9170 ;
      RECT 0.2790 0.6320 0.9370 0.6480 ;
      RECT 0.8870 0.2730 0.9370 0.5820 ;
      RECT 0.2790 0.2760 0.3290 0.5980 ;
      RECT 0.7350 1.0180 1.0890 1.0680 ;
      RECT 1.0390 1.0680 1.0890 1.5680 ;
      RECT 0.7350 1.0680 0.7850 1.2230 ;
      RECT 0.5830 1.3230 0.6330 1.5500 ;
      RECT 0.8870 1.3230 0.9370 1.5570 ;
      RECT 0.2790 1.2730 0.9370 1.3230 ;
      RECT 0.2790 1.3230 0.3290 1.5570 ;
    LAYER PO ;
      RECT 1.7330 0.0700 1.7630 1.6110 ;
      RECT 1.2770 0.0750 1.3070 1.6160 ;
      RECT 1.4290 0.0780 1.4590 1.6180 ;
      RECT 1.5810 0.0660 1.6110 1.6180 ;
      RECT 1.8850 0.0700 1.9150 1.6110 ;
      RECT 0.6690 0.0720 0.6990 1.6210 ;
      RECT 0.5170 0.0720 0.5470 1.6210 ;
      RECT 0.3650 0.0670 0.3950 1.6210 ;
      RECT 0.0610 0.0720 0.0910 1.6210 ;
      RECT 0.9730 0.0760 1.0030 1.6210 ;
      RECT 0.8210 0.0720 0.8510 1.6210 ;
      RECT 0.2130 0.0720 0.2430 1.6210 ;
      RECT 1.1250 0.0760 1.1550 1.6210 ;
  END
END AO221X2_LVT

MACRO AO222X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.976 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1590 0.2490 1.2710 0.3590 ;
        RECT 1.1590 0.3590 1.2090 0.5390 ;
        RECT 1.1590 0.5390 1.3330 0.5890 ;
    END
    ANTENNAGATEAREA 0.0249 ;
  END A6

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7030 0.0970 0.8630 0.2070 ;
    END
    ANTENNAGATEAREA 0.0249 ;
  END A3

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.9760 0.0300 ;
        RECT 1.4950 0.0300 1.5450 0.4840 ;
        RECT 0.5830 0.0300 0.6330 0.4800 ;
        RECT 1.3430 0.0300 1.3930 0.4660 ;
    END
  END VSS

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3990 0.5530 0.5560 0.6630 ;
    END
    ANTENNAGATEAREA 0.0249 ;
  END A2

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.9760 1.7020 ;
        RECT 1.4950 1.0120 1.5450 1.6420 ;
        RECT 0.4310 1.3730 0.4810 1.6420 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6170 1.1610 1.7270 1.2710 ;
        RECT 1.6470 1.2710 1.6970 1.5540 ;
        RECT 1.6470 0.8640 1.6970 1.1610 ;
        RECT 1.6470 0.8030 1.7470 0.8640 ;
        RECT 1.6970 0.4840 1.7470 0.8030 ;
        RECT 1.6470 0.4340 1.7470 0.4840 ;
        RECT 1.6470 0.1260 1.6970 0.4340 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.0090 0.6630 1.1190 ;
        RECT 0.6120 0.8890 0.6620 1.0090 ;
        RECT 0.6120 0.8390 0.7250 0.8890 ;
    END
    ANTENNAGATEAREA 0.0249 ;
  END A4

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2470 0.8570 0.4050 0.9670 ;
        RECT 0.3550 0.8250 0.4050 0.8570 ;
    END
    ANTENNAGATEAREA 0.0249 ;
  END A1

  PIN A5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0070 0.7050 1.1170 0.7590 ;
        RECT 1.0070 0.7590 1.1810 0.8090 ;
        RECT 1.0070 0.8090 1.1170 0.8150 ;
    END
    ANTENNAGATEAREA 0.0249 ;
  END A5
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 2.0910 1.7730 ;
    LAYER M1 ;
      RECT 1.4610 0.6360 1.6370 0.6860 ;
      RECT 1.4610 0.6860 1.5110 0.9070 ;
      RECT 1.1900 0.9070 1.5110 0.9080 ;
      RECT 0.8870 0.9080 1.5110 0.9570 ;
      RECT 1.1900 0.8940 1.2400 0.9070 ;
      RECT 0.8870 0.9570 1.2400 0.9580 ;
      RECT 1.1900 0.9580 1.2400 1.4700 ;
      RECT 0.8870 0.3130 1.0890 0.3630 ;
      RECT 1.0390 0.3630 1.0890 0.4870 ;
      RECT 0.8870 0.7670 0.9370 0.9080 ;
      RECT 0.2790 0.7170 0.9370 0.7670 ;
      RECT 0.8870 0.3630 0.9370 0.7170 ;
      RECT 0.2790 0.3180 0.3290 0.7170 ;
      RECT 1.3420 1.1720 1.3920 1.5340 ;
      RECT 1.0390 1.5340 1.3920 1.5840 ;
      RECT 1.0390 1.0710 1.0890 1.5340 ;
      RECT 0.7350 1.0210 1.0890 1.0710 ;
      RECT 0.7350 1.0710 0.7850 1.2230 ;
      RECT 0.7350 1.0110 0.7850 1.0210 ;
      RECT 0.5830 1.3230 0.6330 1.5570 ;
      RECT 0.8870 1.3230 0.9370 1.5570 ;
      RECT 0.2790 1.2730 0.9370 1.3230 ;
      RECT 0.2790 1.3230 0.3290 1.5570 ;
    LAYER PO ;
      RECT 1.7330 0.0750 1.7630 1.6160 ;
      RECT 1.4290 0.0750 1.4590 1.6160 ;
      RECT 1.2770 0.0760 1.3070 1.6210 ;
      RECT 0.6690 0.0720 0.6990 1.6210 ;
      RECT 0.5170 0.0720 0.5470 1.6210 ;
      RECT 0.3650 0.0670 0.3950 1.6210 ;
      RECT 1.8850 0.0750 1.9150 1.6160 ;
      RECT 0.0610 0.0720 0.0910 1.6210 ;
      RECT 0.9730 0.0760 1.0030 1.6210 ;
      RECT 1.5810 0.0760 1.6110 1.6160 ;
      RECT 0.8210 0.0720 0.8510 1.6210 ;
      RECT 0.2130 0.0720 0.2430 1.6210 ;
      RECT 1.1250 0.0760 1.1550 1.6210 ;
  END
END AO222X1_LVT

MACRO AO222X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.128 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0090 0.6990 1.1190 0.7210 ;
        RECT 1.0090 0.7210 1.1810 0.7710 ;
        RECT 1.0090 0.7710 1.1190 0.8150 ;
    END
    ANTENNAGATEAREA 0.03 ;
  END A5

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3550 0.7050 0.4050 0.8570 ;
        RECT 0.2490 0.8570 0.4050 0.9670 ;
    END
    ANTENNAGATEAREA 0.03 ;
  END A1

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.0090 0.6630 1.1190 ;
        RECT 0.6130 0.7600 0.6630 1.0090 ;
        RECT 0.6130 0.7100 0.7250 0.7600 ;
    END
    ANTENNAGATEAREA 0.03 ;
  END A4

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.1280 1.7020 ;
        RECT 1.6470 1.2650 1.6970 1.6420 ;
        RECT 0.4310 1.3730 0.4810 1.6420 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7690 1.0090 1.8790 1.1190 ;
        RECT 1.8000 1.1190 1.8500 1.4700 ;
        RECT 1.8000 0.7830 1.8500 1.0090 ;
        RECT 1.8000 0.7290 1.8880 0.7830 ;
        RECT 1.8380 0.5530 1.8880 0.7290 ;
        RECT 1.4710 0.5030 1.8880 0.5530 ;
        RECT 1.8000 0.4820 1.8880 0.5030 ;
        RECT 1.4710 0.5530 1.5210 0.7440 ;
        RECT 1.4950 0.1740 1.5450 0.5030 ;
        RECT 1.8000 0.1740 1.8500 0.4820 ;
        RECT 1.4710 0.7440 1.5450 0.8060 ;
        RECT 1.4950 0.8060 1.5450 1.1020 ;
    END
    ANTENNADIFFAREA 0.2484 ;
  END Y

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4910 0.4950 0.8160 0.5450 ;
        RECT 0.7050 0.4010 0.8150 0.4950 ;
    END
    ANTENNAGATEAREA 0.03 ;
  END A2

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.1280 0.0300 ;
        RECT 1.3430 0.0300 1.3930 0.4570 ;
        RECT 1.6470 0.0300 1.6970 0.3940 ;
        RECT 0.5830 0.0300 0.6330 0.4390 ;
    END
  END VSS

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 0.0970 0.8150 0.1020 ;
        RECT 0.7050 0.1020 0.8770 0.1520 ;
        RECT 0.7050 0.1520 0.8150 0.2070 ;
    END
    ANTENNAGATEAREA 0.03 ;
  END A3

  PIN A6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 0.4010 1.2840 0.5110 ;
        RECT 1.2340 0.5110 1.2840 0.5130 ;
        RECT 1.2340 0.5130 1.3330 0.5630 ;
    END
    ANTENNAGATEAREA 0.03 ;
  END A6
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 2.2430 1.7730 ;
    LAYER M1 ;
      RECT 1.5710 0.6030 1.7730 0.6790 ;
      RECT 1.5710 0.6790 1.7500 0.6850 ;
      RECT 1.6450 0.6850 1.6950 1.1520 ;
      RECT 1.6450 1.2020 1.6950 1.2050 ;
      RECT 1.1900 1.1520 1.6950 1.2020 ;
      RECT 1.1900 1.2020 1.2400 1.4700 ;
      RECT 1.1900 0.9710 1.2400 1.1520 ;
      RECT 0.8870 0.9210 1.2400 0.9710 ;
      RECT 1.1900 0.9070 1.2400 0.9210 ;
      RECT 0.2790 0.2800 0.3290 0.5970 ;
      RECT 0.8870 0.2890 1.0890 0.3390 ;
      RECT 1.0390 0.3390 1.0890 0.4630 ;
      RECT 0.8870 0.6470 0.9370 0.9210 ;
      RECT 0.2790 0.5970 0.9390 0.6470 ;
      RECT 0.8870 0.3390 0.9370 0.5970 ;
      RECT 0.7350 1.0210 1.0890 1.0710 ;
      RECT 1.0390 1.0710 1.0890 1.5200 ;
      RECT 0.7350 1.0710 0.7850 1.2230 ;
      RECT 1.0390 1.5200 1.3930 1.5700 ;
      RECT 1.3430 1.2860 1.3930 1.5200 ;
      RECT 0.8870 1.3230 0.9370 1.5570 ;
      RECT 0.5830 1.3230 0.6330 1.5570 ;
      RECT 0.2790 1.2730 0.9370 1.3230 ;
      RECT 0.2790 1.3230 0.3290 1.5570 ;
    LAYER PO ;
      RECT 1.4290 0.0750 1.4590 1.6160 ;
      RECT 1.8850 0.0750 1.9150 1.6160 ;
      RECT 1.1250 0.0760 1.1550 1.6210 ;
      RECT 0.2130 0.0720 0.2430 1.6210 ;
      RECT 0.8210 0.0720 0.8510 1.6210 ;
      RECT 1.7330 0.0660 1.7630 1.6180 ;
      RECT 0.9730 0.0760 1.0030 1.6210 ;
      RECT 1.5810 0.0780 1.6110 1.6180 ;
      RECT 0.0610 0.0720 0.0910 1.6210 ;
      RECT 2.0370 0.0750 2.0670 1.6160 ;
      RECT 0.3650 0.0670 0.3950 1.6210 ;
      RECT 0.5170 0.0720 0.5470 1.6210 ;
      RECT 0.6690 0.0720 0.6990 1.6210 ;
      RECT 1.2770 0.0760 1.3070 1.6210 ;
  END
END AO222X2_LVT

MACRO AO22X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.52 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5070 0.9200 0.5570 1.0090 ;
        RECT 0.4010 1.0090 0.5570 1.1190 ;
    END
    ANTENNAGATEAREA 0.0234 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 0.0880 0.8630 0.2170 ;
    END
    ANTENNAGATEAREA 0.0234 ;
  END A3

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.5200 0.0300 ;
        RECT 1.0390 0.0300 1.0890 0.5030 ;
        RECT 0.5830 0.0300 0.6330 0.4020 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.5200 1.7020 ;
        RECT 1.0390 0.8400 1.0890 1.6420 ;
        RECT 0.4310 1.3580 0.4810 1.6420 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.1610 1.2710 1.2710 ;
        RECT 1.1910 1.2710 1.2410 1.5370 ;
        RECT 1.1910 0.8360 1.2410 1.1610 ;
        RECT 1.1910 0.7860 1.2810 0.8360 ;
        RECT 1.2310 0.5040 1.2810 0.7860 ;
        RECT 1.1910 0.4380 1.2810 0.5040 ;
        RECT 1.1910 0.1450 1.2410 0.4380 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 0.5530 0.7080 0.6630 ;
    END
    ANTENNAGATEAREA 0.0234 ;
  END A4

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7050 0.4040 0.8150 ;
    END
    ANTENNAGATEAREA 0.0234 ;
  END A1
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.6350 1.7730 ;
    LAYER M1 ;
      RECT 0.7350 0.8130 0.8080 0.8630 ;
      RECT 0.7350 0.8630 0.7850 1.2080 ;
      RECT 0.8870 0.5030 0.9370 0.5680 ;
      RECT 0.8870 0.3010 0.9370 0.4530 ;
      RECT 0.7580 0.6180 1.1810 0.6680 ;
      RECT 0.7580 0.6680 0.8080 0.8130 ;
      RECT 0.7580 0.5030 0.8080 0.6180 ;
      RECT 0.2790 0.4530 0.9370 0.5030 ;
      RECT 0.2790 0.5030 0.3290 0.5700 ;
      RECT 0.2790 0.3040 0.3290 0.4530 ;
      RECT 0.5830 1.3080 0.6330 1.5430 ;
      RECT 0.8870 1.3080 0.9370 1.5420 ;
      RECT 0.2790 1.2580 0.9370 1.3080 ;
      RECT 0.2790 1.3080 0.3290 1.5420 ;
    LAYER PO ;
      RECT 1.2770 0.0750 1.3070 1.6160 ;
      RECT 0.6690 0.0720 0.6990 1.6210 ;
      RECT 0.5170 0.0720 0.5470 1.6210 ;
      RECT 0.3650 0.0670 0.3950 1.6210 ;
      RECT 1.4290 0.0750 1.4590 1.6160 ;
      RECT 0.0610 0.0720 0.0910 1.6210 ;
      RECT 0.9730 0.0760 1.0030 1.6210 ;
      RECT 1.1250 0.0760 1.1550 1.6160 ;
      RECT 0.8210 0.0720 0.8510 1.6210 ;
      RECT 0.2130 0.0720 0.2430 1.6210 ;
  END
END AO22X1_LVT

MACRO AO22X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.672 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3130 0.7100 1.4320 0.8200 ;
        RECT 1.3440 0.8200 1.3940 1.4700 ;
        RECT 1.3820 0.5180 1.4320 0.7100 ;
        RECT 1.3440 0.4680 1.4320 0.5180 ;
        RECT 1.3440 0.3940 1.3940 0.4680 ;
        RECT 1.0390 0.3440 1.3940 0.3940 ;
        RECT 1.0390 0.1600 1.0890 0.3440 ;
        RECT 1.3440 0.1600 1.3940 0.3440 ;
        RECT 1.0390 0.3940 1.0890 0.4680 ;
        RECT 1.0110 0.4680 1.0890 0.5180 ;
        RECT 1.0110 0.5180 1.0610 0.7300 ;
        RECT 1.0110 0.7300 1.0890 0.7920 ;
        RECT 1.0390 0.7920 1.0890 1.0880 ;
    END
    ANTENNADIFFAREA 0.2484 ;
  END Y

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 0.5530 0.7080 0.6630 ;
    END
    ANTENNAGATEAREA 0.0246 ;
  END A4

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.6720 1.7020 ;
        RECT 0.4310 1.3730 0.4810 1.6420 ;
        RECT 1.1910 1.2510 1.2410 1.6420 ;
    END
  END VDD

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5070 0.8660 0.5570 1.0080 ;
        RECT 0.4010 1.0080 0.5570 1.1180 ;
    END
    ANTENNAGATEAREA 0.0246 ;
  END A2

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.6720 0.0300 ;
        RECT 1.1910 0.0300 1.2410 0.2930 ;
        RECT 0.5830 0.0300 0.6330 0.4030 ;
    END
  END VSS

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7050 0.4040 0.8150 ;
    END
    ANTENNAGATEAREA 0.0246 ;
  END A1

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 0.0970 0.8630 0.2070 ;
    END
    ANTENNAGATEAREA 0.0246 ;
  END A3
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.7870 1.7730 ;
    LAYER M1 ;
      RECT 1.1150 0.5740 1.3170 0.6560 ;
      RECT 1.1890 0.6560 1.2390 1.1380 ;
      RECT 0.7350 1.1380 1.2390 1.1880 ;
      RECT 0.2790 0.5030 0.3290 0.5360 ;
      RECT 0.2790 0.2700 0.3290 0.4530 ;
      RECT 0.7350 1.1880 0.7850 1.1890 ;
      RECT 0.7350 1.0150 0.7850 1.1380 ;
      RECT 0.8870 0.5030 0.9370 1.1380 ;
      RECT 0.8870 0.2700 0.9370 0.4530 ;
      RECT 0.2790 0.4530 0.9370 0.5030 ;
      RECT 0.8870 1.3230 0.9370 1.5570 ;
      RECT 0.5830 1.3230 0.6330 1.5570 ;
      RECT 0.2790 1.2730 0.9370 1.3230 ;
      RECT 0.2790 1.3230 0.3290 1.5570 ;
    LAYER PO ;
      RECT 1.4290 0.0560 1.4590 1.5970 ;
      RECT 1.2770 0.0520 1.3070 1.6040 ;
      RECT 1.5810 0.0560 1.6110 1.5970 ;
      RECT 1.1250 0.0640 1.1550 1.6040 ;
      RECT 0.2130 0.0720 0.2430 1.6210 ;
      RECT 0.8210 0.0720 0.8510 1.6210 ;
      RECT 0.9730 0.0760 1.0030 1.6210 ;
      RECT 0.0610 0.0720 0.0910 1.6210 ;
      RECT 0.3650 0.0670 0.3950 1.6210 ;
      RECT 0.5170 0.0720 0.5470 1.6210 ;
      RECT 0.6690 0.0720 0.6990 1.6210 ;
  END
END AO22X2_LVT

MACRO AOBUFX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.28 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1570 0.7470 1.3330 0.8070 ;
        RECT 1.1610 0.8070 1.2710 0.8150 ;
        RECT 1.1610 0.7050 1.2710 0.7470 ;
    END
    ANTENNAGATEAREA 0.0306 ;
  END A

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.8180 1.0090 1.0080 1.1190 ;
        RECT 0.8820 0.9910 0.9420 1.0090 ;
        RECT 0.8820 1.1190 0.9420 1.2870 ;
        RECT 0.8820 1.2870 1.2410 1.3370 ;
        RECT 1.1910 1.3370 1.2410 1.4280 ;
        RECT 1.1910 0.8860 1.2410 1.2870 ;
    END
  END VDDG

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.2800 1.7020 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0460 2.5130 1.2410 2.5630 ;
        RECT 1.1910 1.9290 1.2410 2.5130 ;
        RECT 1.0460 2.5630 1.0960 2.6810 ;
        RECT 1.0090 2.6810 1.1190 2.7570 ;
        RECT 1.0090 2.7570 1.2410 2.8070 ;
        RECT 1.1910 2.8070 1.2410 3.1550 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.2800 0.0300 ;
        RECT 1.1910 0.0300 1.2410 0.6140 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 2.2800 3.3740 ;
        RECT 1.3430 2.7820 1.3930 3.3140 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT 0.7930 0.6790 1.6180 2.6650 ;
    LAYER M1 ;
      RECT 0.9470 1.8100 1.3930 1.8600 ;
      RECT 1.3430 1.8600 1.3930 2.5640 ;
      RECT 1.2510 2.6140 1.6370 2.6740 ;
      RECT 1.3270 1.1760 1.5380 1.2260 ;
      RECT 1.3430 1.2260 1.3930 1.4280 ;
      RECT 1.4880 0.5610 1.5380 1.1760 ;
      RECT 1.3430 0.5110 1.6370 0.5610 ;
      RECT 1.3430 0.5610 1.3930 0.6140 ;
      RECT 1.3430 0.2560 1.3930 0.5110 ;
    LAYER PO ;
      RECT 2.0370 0.1330 2.0670 1.4920 ;
      RECT 2.0370 1.7230 2.0670 3.2150 ;
      RECT 0.0610 1.7230 0.0910 3.2150 ;
      RECT 0.0610 0.1340 0.0910 1.4930 ;
      RECT 2.1890 1.7230 2.2190 3.2150 ;
      RECT 2.1890 0.1330 2.2190 1.4920 ;
      RECT 1.1250 1.7230 1.1550 3.2150 ;
      RECT 1.5810 0.1340 1.6110 3.2150 ;
      RECT 0.8210 1.7230 0.8510 3.2150 ;
      RECT 0.8210 0.1340 0.8510 1.4980 ;
      RECT 0.9730 0.1340 1.0030 3.2150 ;
      RECT 1.8850 1.7230 1.9150 3.2150 ;
      RECT 1.7330 1.7230 1.7630 3.2150 ;
      RECT 0.6690 1.7230 0.6990 3.2150 ;
      RECT 1.2770 1.7230 1.3070 3.2150 ;
      RECT 0.5170 1.7230 0.5470 3.2150 ;
      RECT 0.3650 1.7230 0.3950 3.2150 ;
      RECT 0.2130 1.7230 0.2430 3.2150 ;
      RECT 1.4290 1.7230 1.4590 3.2150 ;
      RECT 0.6690 0.1340 0.6990 1.4930 ;
      RECT 0.5170 0.1340 0.5470 1.4930 ;
      RECT 0.3650 0.1340 0.3950 1.4930 ;
      RECT 0.2130 0.1340 0.2430 1.4930 ;
      RECT 1.7330 0.1330 1.7630 1.4920 ;
      RECT 1.8850 0.1330 1.9150 1.4920 ;
      RECT 1.1250 0.1340 1.1550 1.4980 ;
      RECT 1.2770 0.1340 1.3070 1.4980 ;
      RECT 1.4290 0.1340 1.4590 1.4980 ;
  END
END AOBUFX1_LVT

MACRO AOBUFX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.432 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 0.7660 1.3330 0.8260 ;
        RECT 1.1610 0.7060 1.2710 0.7660 ;
    END
    ANTENNAGATEAREA 0.0306 ;
  END A

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.8180 1.0090 1.0080 1.1190 ;
        RECT 0.8820 0.9910 0.9420 1.0090 ;
        RECT 0.8820 1.1190 0.9420 1.3060 ;
        RECT 0.8820 1.3060 1.2410 1.3560 ;
        RECT 1.1910 1.3560 1.2410 1.4470 ;
        RECT 1.1910 0.9970 1.2410 1.3060 ;
    END
  END VDDG

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.4320 1.7020 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0460 2.5040 1.5450 2.5540 ;
        RECT 1.1910 1.9200 1.2410 2.5040 ;
        RECT 1.4950 1.8280 1.5450 2.5040 ;
        RECT 1.0460 2.5540 1.0960 2.6820 ;
        RECT 1.0090 2.6820 1.1190 2.7570 ;
        RECT 1.0090 2.7570 1.5450 2.8070 ;
        RECT 1.0090 2.8070 1.1190 2.8080 ;
        RECT 1.1910 2.8070 1.2410 3.1550 ;
        RECT 1.4950 2.8070 1.5450 3.1550 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END Y

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.4320 0.0300 ;
        RECT 1.1910 0.0300 1.2410 0.5420 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 2.4320 3.3740 ;
        RECT 1.3430 2.8910 1.3930 3.3140 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT 0.7910 0.6790 1.7690 2.6650 ;
    LAYER M1 ;
      RECT 0.9470 1.8100 1.3930 1.8600 ;
      RECT 1.3430 1.8600 1.3930 2.4190 ;
      RECT 1.3430 1.7830 1.3930 1.8100 ;
      RECT 1.2510 2.6140 1.6370 2.6740 ;
      RECT 1.3270 1.1950 1.5380 1.2450 ;
      RECT 1.3430 1.2450 1.3930 1.4470 ;
      RECT 1.3430 0.9010 1.3930 1.1950 ;
      RECT 1.4880 0.4940 1.5380 1.1950 ;
      RECT 1.3430 0.4440 1.6370 0.4940 ;
      RECT 1.3430 0.4940 1.3930 0.6140 ;
      RECT 1.3430 0.2560 1.3930 0.4440 ;
    LAYER PO ;
      RECT 0.3650 1.7230 0.3950 3.2150 ;
      RECT 0.5170 1.7230 0.5470 3.2150 ;
      RECT 0.6690 1.7230 0.6990 3.2150 ;
      RECT 1.8850 1.7230 1.9150 3.2150 ;
      RECT 2.0370 1.7230 2.0670 3.2150 ;
      RECT 2.1890 1.7230 2.2190 3.2150 ;
      RECT 0.2130 1.7230 0.2430 3.2150 ;
      RECT 0.6690 0.1370 0.6990 1.5140 ;
      RECT 0.5170 0.1370 0.5470 1.5140 ;
      RECT 0.3650 0.1370 0.3950 1.5140 ;
      RECT 0.2130 0.1370 0.2430 1.5140 ;
      RECT 2.1890 0.1320 2.2190 1.5170 ;
      RECT 2.0370 0.1320 2.0670 1.5170 ;
      RECT 1.8850 0.1320 1.9150 1.5170 ;
      RECT 0.0610 0.1370 0.0910 1.5140 ;
      RECT 1.1250 1.7230 1.1550 3.2150 ;
      RECT 0.0610 1.7230 0.0910 3.2150 ;
      RECT 2.3410 0.1320 2.3710 1.5170 ;
      RECT 2.3410 1.7230 2.3710 3.2150 ;
      RECT 1.7330 0.1340 1.7630 1.5170 ;
      RECT 1.7330 1.7230 1.7630 3.2150 ;
      RECT 1.5810 0.1340 1.6110 3.2150 ;
      RECT 0.8210 1.7230 0.8510 3.2150 ;
      RECT 0.8210 0.1340 0.8510 1.5170 ;
      RECT 0.9730 0.1340 1.0030 3.2150 ;
      RECT 1.2770 1.7230 1.3070 3.2150 ;
      RECT 1.4290 1.7230 1.4590 3.2150 ;
      RECT 1.1250 0.1340 1.1550 1.5170 ;
      RECT 1.2770 0.1340 1.3070 1.5170 ;
      RECT 1.4290 0.1340 1.4590 1.5170 ;
  END
END AOBUFX2_LVT

MACRO AOBUFX4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.432 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0090 0.8690 1.1810 0.9290 ;
        RECT 1.0090 0.8570 1.1190 0.8690 ;
        RECT 1.0090 0.9290 1.1190 0.9670 ;
    END
    ANTENNAGATEAREA 0.0306 ;
  END A

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.6660 1.0090 0.8560 1.1190 ;
        RECT 0.7300 0.9910 0.7900 1.0090 ;
        RECT 0.7300 1.1190 0.7900 1.4200 ;
        RECT 0.7300 1.4200 1.0890 1.4700 ;
        RECT 1.0390 1.4700 1.0890 1.5600 ;
        RECT 1.0390 1.0180 1.0890 1.4200 ;
    END
  END VDDG

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.4320 1.7020 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8940 2.5040 1.6970 2.5540 ;
        RECT 1.0390 1.9200 1.0890 2.5040 ;
        RECT 1.3430 1.9200 1.3930 2.5040 ;
        RECT 1.6470 1.9200 1.6970 2.5040 ;
        RECT 0.8940 2.5540 0.9440 2.6810 ;
        RECT 0.8570 2.6810 0.9670 2.7570 ;
        RECT 0.8570 2.7570 1.6970 2.8070 ;
        RECT 1.6470 2.8070 1.6970 3.1550 ;
        RECT 1.0390 2.8070 1.0890 3.1550 ;
        RECT 1.3430 2.8070 1.3930 3.1550 ;
    END
    ANTENNADIFFAREA 0.3976 ;
  END Y

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.4320 0.0300 ;
        RECT 1.0390 0.0300 1.0890 0.5420 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 2.4320 3.3740 ;
        RECT 1.4950 2.8910 1.5450 3.3140 ;
        RECT 1.1910 2.8910 1.2410 3.3140 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT 0.6420 0.6790 1.7780 2.6650 ;
    LAYER M1 ;
      RECT 0.7950 1.8100 1.5450 1.8600 ;
      RECT 1.4950 1.8600 1.5450 2.4190 ;
      RECT 1.4950 1.7830 1.5450 1.8100 ;
      RECT 1.1910 1.8600 1.2410 2.4190 ;
      RECT 1.1910 1.7830 1.2410 1.8100 ;
      RECT 1.0990 2.6140 1.6370 2.6740 ;
      RECT 1.1910 1.3080 1.3860 1.3580 ;
      RECT 1.1910 1.3580 1.2410 1.5600 ;
      RECT 1.1910 1.0140 1.2410 1.3080 ;
      RECT 1.3360 1.3580 1.3860 1.3590 ;
      RECT 1.3360 0.5870 1.3860 1.3080 ;
      RECT 1.1910 0.5370 1.4850 0.5870 ;
      RECT 1.1910 0.5870 1.2410 0.6140 ;
      RECT 1.1910 0.2560 1.2410 0.5370 ;
    LAYER PO ;
      RECT 2.3410 1.7230 2.3710 3.2150 ;
      RECT 2.1890 1.7230 2.2190 3.2150 ;
      RECT 2.0370 1.7230 2.0670 3.2150 ;
      RECT 1.8850 1.7230 1.9150 3.2150 ;
      RECT 0.5170 1.7230 0.5470 3.2150 ;
      RECT 0.3650 1.7230 0.3950 3.2150 ;
      RECT 1.5810 1.7230 1.6110 3.2150 ;
      RECT 1.5810 0.1330 1.6110 1.6230 ;
      RECT 0.9730 1.7230 1.0030 3.2150 ;
      RECT 1.7330 0.1330 1.7630 1.6230 ;
      RECT 1.7330 1.7230 1.7630 3.2150 ;
      RECT 0.2130 1.7230 0.2430 3.2150 ;
      RECT 0.0610 1.7230 0.0910 3.2150 ;
      RECT 1.4290 0.1340 1.4590 3.2150 ;
      RECT 0.6690 1.7230 0.6990 3.2150 ;
      RECT 0.6690 0.1340 0.6990 1.6230 ;
      RECT 0.8210 0.1340 0.8510 3.2150 ;
      RECT 2.1890 0.1330 2.2190 1.6230 ;
      RECT 2.0370 0.1330 2.0670 1.6230 ;
      RECT 1.8850 0.1330 1.9150 1.6230 ;
      RECT 1.1250 1.7230 1.1550 3.2150 ;
      RECT 1.2770 1.7230 1.3070 3.2150 ;
      RECT 0.5170 0.1330 0.5470 1.6230 ;
      RECT 0.3650 0.1330 0.3950 1.6230 ;
      RECT 0.2130 0.1330 0.2430 1.6230 ;
      RECT 0.9730 0.1330 1.0030 1.6230 ;
      RECT 1.1250 0.1330 1.1550 1.6230 ;
      RECT 0.0610 0.1330 0.0910 1.6230 ;
      RECT 1.2770 0.1330 1.3070 1.6230 ;
      RECT 2.3410 0.1330 2.3710 1.6230 ;
  END
END AOBUFX4_LVT

MACRO AODFFARX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.584 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 2.3770 0.3590 2.4370 ;
        RECT 0.2490 2.4370 0.6330 2.4870 ;
        RECT 0.2490 2.4870 0.2990 3.0110 ;
        RECT 0.5830 1.8950 0.6330 2.4370 ;
        RECT 0.2490 3.0110 0.6330 3.0610 ;
        RECT 0.5830 3.0610 0.6330 3.2220 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.4620 0.7250 1.5910 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6970 0.3590 0.7020 ;
        RECT 0.2490 0.7020 0.4210 0.7520 ;
        RECT 0.2490 0.7520 0.3590 0.8140 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7230 0.1580 1.8790 0.2070 ;
        RECT 1.7230 0.1080 2.5490 0.1580 ;
        RECT 1.7230 0.0970 1.8790 0.1080 ;
    END
    ANTENNAGATEAREA 0.0441 ;
  END RSTB

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0970 2.1230 0.2070 2.1830 ;
        RECT 0.0970 2.0730 0.3290 2.1230 ;
        RECT 0.0970 2.1830 0.1470 3.1420 ;
        RECT 0.2790 1.8950 0.3290 2.0730 ;
        RECT 0.0970 3.1420 0.3450 3.1920 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.2740 1.4230 0.3340 1.5660 ;
        RECT 0.2210 1.3380 0.3760 1.4230 ;
        RECT 0.0350 1.2880 0.9370 1.3380 ;
        RECT 0.8870 1.3380 0.9370 1.3910 ;
        RECT 0.2740 1.0550 0.3340 1.2880 ;
        RECT 0.7350 1.1200 0.7850 1.2880 ;
        RECT 0.7350 1.3380 0.7850 1.3860 ;
        RECT 0.8870 1.1330 0.9370 1.2880 ;
        RECT 0.8870 1.3910 2.0170 1.4410 ;
    END
  END VDDG

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.5840 1.7020 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.5840 0.0300 ;
        RECT 0.5860 0.0300 0.6360 0.2180 ;
        RECT 0.2790 0.0300 0.3290 0.4410 ;
        RECT 1.5410 0.0300 1.5910 0.3090 ;
        RECT 0.5860 0.2180 0.9370 0.2680 ;
        RECT 1.5410 0.3090 2.0010 0.3590 ;
        RECT 0.7350 0.2680 0.7850 0.4720 ;
        RECT 0.8870 0.2680 0.9370 0.4720 ;
        RECT 1.9510 0.3590 2.0010 0.4830 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 2.5840 3.3740 ;
        RECT 0.4310 3.1340 0.4810 3.3140 ;
        RECT 1.0150 3.0490 1.0650 3.3140 ;
        RECT 1.0150 2.9990 2.1690 3.0490 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 2.6990 2.6650 ;
    LAYER M1 ;
      RECT 0.6950 2.1120 0.8200 2.1620 ;
      RECT 0.6950 2.1620 0.7450 2.5710 ;
      RECT 0.3550 2.5710 0.7450 2.6210 ;
      RECT 0.3550 2.8820 1.6970 2.9320 ;
      RECT 1.3440 2.6040 1.3940 2.8820 ;
      RECT 1.6470 2.6010 1.6970 2.8820 ;
      RECT 1.2510 2.5540 1.3940 2.6040 ;
      RECT 1.6070 2.5510 1.6970 2.6010 ;
      RECT 1.6070 2.3640 1.6570 2.5510 ;
      RECT 1.6070 2.3140 1.7150 2.3640 ;
      RECT 0.3550 2.6210 0.4050 2.8820 ;
      RECT 1.1750 0.3370 1.2650 0.3870 ;
      RECT 1.2150 0.3870 1.2650 1.0100 ;
      RECT 0.4310 1.0100 1.2650 1.0600 ;
      RECT 1.1910 1.0600 1.2410 1.3360 ;
      RECT 0.4310 0.8510 0.4810 1.0100 ;
      RECT 0.4310 0.6010 0.5210 0.6510 ;
      RECT 0.4310 0.4770 0.4810 0.6010 ;
      RECT 0.4310 0.8020 0.5210 0.8510 ;
      RECT 0.4710 0.6510 0.5210 0.8020 ;
      RECT 0.4310 1.0600 0.4810 1.2380 ;
      RECT 1.3430 1.1800 2.2450 1.2300 ;
      RECT 1.3430 1.2300 1.3930 1.3360 ;
      RECT 1.3430 1.0720 1.3930 1.1800 ;
      RECT 1.3150 1.0190 1.3930 1.0720 ;
      RECT 1.3150 0.7680 1.3650 1.0190 ;
      RECT 1.3150 0.7100 1.3930 0.7680 ;
      RECT 1.3430 0.5060 1.3930 0.7100 ;
      RECT 1.3430 0.3770 1.3930 0.4560 ;
      RECT 1.3430 0.4560 1.5610 0.5060 ;
      RECT 1.8100 2.6360 1.9510 2.6860 ;
      RECT 1.8100 2.4640 1.8600 2.6360 ;
      RECT 1.7070 2.4140 1.8600 2.4640 ;
      RECT 1.8100 2.2260 1.8600 2.4140 ;
      RECT 0.9630 2.1760 1.8600 2.2260 ;
      RECT 0.9630 2.2260 1.0130 2.6610 ;
      RECT 0.0350 1.7610 2.1290 1.8170 ;
      RECT 0.6950 1.8170 0.7450 2.0120 ;
      RECT 2.0790 1.8170 2.1290 2.0420 ;
      RECT 0.6950 2.0120 1.4220 2.0620 ;
      RECT 2.0790 2.0420 2.1690 2.0920 ;
      RECT 0.4310 1.8170 0.4810 2.3410 ;
      RECT 1.9510 2.5330 2.3970 2.5830 ;
      RECT 2.2990 2.5830 2.3490 2.8950 ;
      RECT 1.9510 2.0620 2.0010 2.5330 ;
      RECT 1.7800 2.8950 2.3490 2.9450 ;
      RECT 1.7820 2.0120 2.0010 2.0620 ;
      RECT 1.0870 1.5400 2.0930 1.5900 ;
      RECT 1.5550 1.0230 2.3970 1.0730 ;
      RECT 1.1150 3.1030 1.9610 3.1530 ;
      RECT 1.1150 3.1530 1.1650 3.2270 ;
      RECT 1.0390 0.5400 1.1650 0.5900 ;
      RECT 1.0390 0.4160 1.0890 0.5400 ;
      RECT 1.1150 0.5900 1.1650 0.7400 ;
      RECT 1.0390 0.7400 1.1650 0.7900 ;
      RECT 1.0390 0.7900 1.0890 0.9360 ;
      RECT 1.4710 2.7740 1.5610 2.8240 ;
      RECT 1.4900 2.4100 1.5400 2.7740 ;
      RECT 1.4900 2.3920 1.5450 2.4100 ;
      RECT 1.1510 2.3420 1.5450 2.3920 ;
      RECT 1.1510 2.3920 1.2010 2.7130 ;
      RECT 1.4950 2.3210 1.5450 2.3420 ;
      RECT 0.4910 2.7130 1.2010 2.7630 ;
      RECT 1.1510 2.7630 1.2010 2.7650 ;
      RECT 0.5830 0.6400 1.0290 0.6900 ;
      RECT 0.5830 0.6900 0.6330 0.9360 ;
      RECT 0.5830 0.4440 0.6330 0.6400 ;
      RECT 1.4030 3.2030 2.5490 3.2530 ;
      RECT 1.4190 0.8590 1.9410 0.9090 ;
      RECT 1.4190 0.9090 1.4690 0.9460 ;
      RECT 2.0110 2.6800 2.2450 2.7300 ;
      RECT 1.8590 0.5620 2.0930 0.6120 ;
      RECT 0.9470 1.8910 1.1820 1.9410 ;
      RECT 0.7810 0.1180 1.4910 0.1680 ;
      RECT 1.4790 1.2860 1.8650 1.3360 ;
    LAYER PO ;
      RECT 0.6690 1.7550 0.6990 3.2820 ;
      RECT 1.7330 2.6520 1.7630 3.2820 ;
      RECT 0.3650 1.7400 0.3950 3.2820 ;
      RECT 1.2770 0.0900 1.3070 0.5640 ;
      RECT 0.8210 1.7550 0.8510 3.2820 ;
      RECT 1.8850 0.7800 1.9150 3.2820 ;
      RECT 0.5170 0.0900 0.5470 1.6280 ;
      RECT 1.5810 0.0900 1.6110 1.6280 ;
      RECT 0.9730 0.0900 1.0030 1.6280 ;
      RECT 1.4290 0.0900 1.4590 1.6280 ;
      RECT 0.8210 0.0900 0.8510 1.6280 ;
      RECT 1.7330 0.0900 1.7630 1.6280 ;
      RECT 0.6690 0.0900 0.6990 1.6280 ;
      RECT 2.0370 0.0900 2.0670 1.6280 ;
      RECT 1.1250 0.0900 1.1550 3.2820 ;
      RECT 0.3650 0.0900 0.3950 1.6280 ;
      RECT 1.5810 1.7550 1.6110 3.2820 ;
      RECT 1.4290 1.7550 1.4590 3.2820 ;
      RECT 0.5170 1.7400 0.5470 3.2820 ;
      RECT 2.0370 1.7550 2.0670 3.2820 ;
      RECT 2.4930 0.0900 2.5230 3.2820 ;
      RECT 1.8850 0.0900 1.9150 0.6400 ;
      RECT 1.2770 1.7550 1.3070 3.2820 ;
      RECT 0.2130 0.2490 0.2430 3.2820 ;
      RECT 2.1890 0.0900 2.2190 3.2820 ;
      RECT 0.9730 2.5610 1.0030 3.2820 ;
      RECT 0.0610 0.2490 0.0910 3.2820 ;
      RECT 2.3410 0.0900 2.3710 3.2820 ;
      RECT 0.9730 1.7550 1.0030 2.3580 ;
      RECT 1.2770 1.0120 1.3070 1.6280 ;
      RECT 1.7330 1.7550 1.7630 2.4920 ;
  END
END AODFFARX1_LVT

MACRO AODFFARX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.888 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 1.4580 1.0290 1.5870 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 0.6970 0.6630 0.7020 ;
        RECT 0.5530 0.7020 0.7250 0.7520 ;
        RECT 0.5530 0.7520 0.6630 0.8140 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0270 0.1080 2.8530 0.1580 ;
        RECT 2.0270 0.0970 2.1830 0.1080 ;
        RECT 2.0270 0.1580 2.1830 0.2070 ;
    END
    ANTENNAGATEAREA 0.0441 ;
  END RSTB

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0970 3.1370 0.2070 3.2470 ;
        RECT 0.1150 3.0800 0.1650 3.1370 ;
        RECT 0.1150 3.0300 0.4810 3.0800 ;
        RECT 0.1150 2.4320 0.1650 3.0300 ;
        RECT 0.4310 3.0800 0.4810 3.2020 ;
        RECT 0.1150 2.3820 0.4810 2.4320 ;
        RECT 0.4310 1.8780 0.4810 2.3820 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2390 2.4960 0.7850 2.5460 ;
        RECT 0.7350 1.8880 0.7850 2.4960 ;
        RECT 0.2390 2.5460 0.2890 2.8330 ;
        RECT 0.2390 2.8330 0.3590 2.9200 ;
        RECT 0.2390 2.9200 0.7850 2.9700 ;
        RECT 0.7350 2.9700 0.7850 3.2020 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.5780 1.4230 0.6380 1.5660 ;
        RECT 0.5250 1.3380 0.6800 1.4230 ;
        RECT 0.0350 1.2880 1.2410 1.3380 ;
        RECT 1.1910 1.3380 1.2410 1.3910 ;
        RECT 0.5780 1.0550 0.6380 1.2880 ;
        RECT 1.0390 1.3380 1.0890 1.3860 ;
        RECT 1.0390 1.1200 1.0890 1.2880 ;
        RECT 1.1910 1.1330 1.2410 1.2880 ;
        RECT 1.1910 1.3910 2.3210 1.4410 ;
    END
  END VDDG

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.8880 1.7020 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.8880 0.0300 ;
        RECT 0.8900 0.0300 0.9400 0.2180 ;
        RECT 0.5830 0.0300 0.6330 0.4410 ;
        RECT 1.8450 0.0300 1.8950 0.3090 ;
        RECT 0.8900 0.2180 1.2410 0.2680 ;
        RECT 1.8450 0.3090 2.3050 0.3590 ;
        RECT 1.0390 0.2680 1.0890 0.4720 ;
        RECT 1.1910 0.2680 1.2410 0.4720 ;
        RECT 2.2550 0.3590 2.3050 0.4830 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 2.8880 3.3740 ;
        RECT 0.5830 3.0380 0.6330 3.3140 ;
        RECT 0.2790 3.1300 0.3290 3.3140 ;
        RECT 0.8870 2.9270 0.9370 3.3140 ;
        RECT 1.3190 3.0490 1.3690 3.3140 ;
        RECT 1.3190 2.9990 2.4730 3.0490 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 3.0030 2.6650 ;
    LAYER M1 ;
      RECT 1.6480 2.8820 2.0010 2.9320 ;
      RECT 1.6480 2.8460 1.6980 2.8820 ;
      RECT 1.9510 2.6010 2.0010 2.8820 ;
      RECT 0.5260 2.7960 1.6980 2.8460 ;
      RECT 1.9110 2.5510 2.0010 2.6010 ;
      RECT 1.6480 2.6040 1.6980 2.7960 ;
      RECT 1.9110 2.3640 1.9610 2.5510 ;
      RECT 1.5550 2.5540 1.6980 2.6040 ;
      RECT 1.9110 2.3140 2.0190 2.3640 ;
      RECT 0.9990 2.1620 1.0490 2.5960 ;
      RECT 0.9990 2.1120 1.1240 2.1620 ;
      RECT 0.5260 2.5960 1.0490 2.6460 ;
      RECT 0.5260 2.8460 0.5760 2.8470 ;
      RECT 0.5260 2.7460 0.5760 2.7960 ;
      RECT 0.3390 2.6960 0.5760 2.7460 ;
      RECT 0.5260 2.6460 0.5760 2.6960 ;
      RECT 1.4790 0.3370 1.5690 0.3870 ;
      RECT 1.5190 0.3870 1.5690 1.0100 ;
      RECT 0.7350 1.0100 1.5690 1.0600 ;
      RECT 1.4950 1.0600 1.5450 1.3360 ;
      RECT 0.7350 0.8510 0.7850 1.0100 ;
      RECT 0.7350 0.6010 0.8250 0.6510 ;
      RECT 0.7350 0.4770 0.7850 0.6010 ;
      RECT 0.7350 0.8020 0.8250 0.8510 ;
      RECT 0.7750 0.6510 0.8250 0.8020 ;
      RECT 0.7350 1.0600 0.7850 1.2380 ;
      RECT 1.6470 1.1800 2.5490 1.2300 ;
      RECT 1.6470 1.2300 1.6970 1.3360 ;
      RECT 1.6470 1.0720 1.6970 1.1800 ;
      RECT 1.6190 1.0190 1.6970 1.0720 ;
      RECT 1.6190 0.7680 1.6690 1.0190 ;
      RECT 1.6190 0.7100 1.6970 0.7680 ;
      RECT 1.6470 0.5060 1.6970 0.7100 ;
      RECT 1.6470 0.3770 1.6970 0.4560 ;
      RECT 1.6470 0.4560 1.8650 0.5060 ;
      RECT 1.4190 3.1040 2.2650 3.1540 ;
      RECT 1.4190 3.1540 1.4690 3.2270 ;
      RECT 1.0850 0.1180 1.7950 0.1680 ;
      RECT 2.3830 2.0420 2.4730 2.0920 ;
      RECT 2.3830 1.8110 2.4330 2.0420 ;
      RECT 0.0350 1.7550 2.4330 1.8110 ;
      RECT 0.8870 1.8110 0.9370 2.4380 ;
      RECT 0.9990 1.8110 1.0490 2.0120 ;
      RECT 0.9990 2.0120 1.7260 2.0620 ;
      RECT 0.5830 1.8110 0.6330 2.3900 ;
      RECT 0.2790 1.8110 0.3290 2.2980 ;
      RECT 2.0860 2.0120 2.3050 2.0620 ;
      RECT 2.2550 2.0620 2.3050 2.5330 ;
      RECT 2.2550 2.5330 2.7010 2.5830 ;
      RECT 2.6030 2.5830 2.6530 2.8950 ;
      RECT 2.0840 2.8950 2.6530 2.9450 ;
      RECT 1.7830 1.2860 2.1690 1.3360 ;
      RECT 2.1140 2.6360 2.2550 2.6860 ;
      RECT 2.1140 2.4640 2.1640 2.6360 ;
      RECT 2.0110 2.4140 2.1640 2.4640 ;
      RECT 2.1140 2.2260 2.1640 2.4140 ;
      RECT 1.2670 2.1760 2.1640 2.2260 ;
      RECT 1.2670 2.2260 1.3170 2.6460 ;
      RECT 1.3910 1.5400 2.3970 1.5900 ;
      RECT 1.8590 1.0230 2.7010 1.0730 ;
      RECT 1.3430 0.5400 1.4690 0.5900 ;
      RECT 1.3430 0.4160 1.3930 0.5400 ;
      RECT 1.4190 0.5900 1.4690 0.7400 ;
      RECT 1.3430 0.7400 1.4690 0.7900 ;
      RECT 1.3430 0.7900 1.3930 0.9360 ;
      RECT 1.7750 2.7740 1.8650 2.8240 ;
      RECT 1.7940 2.4100 1.8440 2.7740 ;
      RECT 1.7940 2.3920 1.8490 2.4100 ;
      RECT 1.4550 2.3420 1.8490 2.3920 ;
      RECT 1.4550 2.3920 1.5050 2.6960 ;
      RECT 1.7990 2.3210 1.8490 2.3420 ;
      RECT 0.6430 2.6960 1.5050 2.7460 ;
      RECT 0.8870 0.6400 1.3330 0.6900 ;
      RECT 0.8870 0.6900 0.9370 0.9360 ;
      RECT 0.8870 0.4440 0.9370 0.6400 ;
      RECT 1.7070 3.2040 2.8530 3.2540 ;
      RECT 1.7230 0.8590 2.2450 0.9090 ;
      RECT 1.7230 0.9090 1.7730 0.9460 ;
      RECT 2.3150 2.6800 2.5490 2.7300 ;
      RECT 2.1630 0.5620 2.3970 0.6120 ;
      RECT 1.2510 1.8910 1.4860 1.9410 ;
    LAYER PO ;
      RECT 0.9730 1.7400 1.0030 3.2820 ;
      RECT 0.8210 1.7400 0.8510 3.2820 ;
      RECT 0.6690 1.7400 0.6990 3.2820 ;
      RECT 0.5170 0.2490 0.5470 3.2820 ;
      RECT 0.0610 0.0900 0.0910 3.2820 ;
      RECT 0.3650 1.7400 0.3950 3.2820 ;
      RECT 0.2130 1.7400 0.2430 3.2820 ;
      RECT 0.2130 0.0900 0.2430 1.6280 ;
      RECT 2.1890 0.0900 2.2190 0.6400 ;
      RECT 1.5810 1.7550 1.6110 3.2820 ;
      RECT 2.4930 0.0900 2.5230 3.2820 ;
      RECT 1.2770 2.5460 1.3070 3.2820 ;
      RECT 2.6450 0.0900 2.6750 3.2820 ;
      RECT 1.2770 1.7550 1.3070 2.3580 ;
      RECT 1.5810 1.0120 1.6110 1.6280 ;
      RECT 2.0370 1.7550 2.0670 2.4920 ;
      RECT 2.0370 2.6520 2.0670 3.2820 ;
      RECT 1.5810 0.0900 1.6110 0.5640 ;
      RECT 1.1250 1.7550 1.1550 3.2820 ;
      RECT 2.1890 0.7800 2.2190 3.2820 ;
      RECT 0.8210 0.0900 0.8510 1.6280 ;
      RECT 1.8850 0.0900 1.9150 1.6280 ;
      RECT 1.2770 0.0900 1.3070 1.6280 ;
      RECT 1.7330 0.0900 1.7630 1.6280 ;
      RECT 1.1250 0.0900 1.1550 1.6280 ;
      RECT 2.0370 0.0900 2.0670 1.6280 ;
      RECT 0.9730 0.0900 1.0030 1.6280 ;
      RECT 2.3410 0.0900 2.3710 1.6280 ;
      RECT 1.4290 0.0900 1.4590 3.2820 ;
      RECT 0.6690 0.0900 0.6990 1.6280 ;
      RECT 1.8850 1.7550 1.9150 3.2820 ;
      RECT 0.3650 0.2490 0.3950 1.6210 ;
      RECT 1.7330 1.7550 1.7630 3.2820 ;
      RECT 2.3410 1.7550 2.3710 3.2820 ;
      RECT 2.7970 0.0900 2.8270 3.2820 ;
  END
END AODFFARX2_LVT

MACRO AODFFNARX1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.584 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 2.3770 0.3590 2.4370 ;
        RECT 0.2490 2.4370 0.6330 2.4870 ;
        RECT 0.2490 2.4870 0.2990 3.0080 ;
        RECT 0.5830 1.8950 0.6330 2.4370 ;
        RECT 0.2490 3.0080 0.6330 3.0580 ;
        RECT 0.2490 3.0580 0.2990 3.0610 ;
        RECT 0.5830 3.0580 0.6330 3.2190 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.4630 0.7250 1.5920 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.6980 0.3590 0.7020 ;
        RECT 0.2490 0.7020 0.4210 0.7520 ;
        RECT 0.2490 0.7520 0.3590 0.8150 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7230 0.1080 2.5490 0.1580 ;
        RECT 1.7230 0.1580 1.8790 0.2070 ;
        RECT 1.7230 0.0970 1.8790 0.1080 ;
    END
    ANTENNAGATEAREA 0.0441 ;
  END RSTB

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0970 2.1230 0.2070 2.1830 ;
        RECT 0.0970 2.0730 0.3290 2.1230 ;
        RECT 0.0970 2.1830 0.1470 3.1630 ;
        RECT 0.2790 1.8950 0.3290 2.0730 ;
        RECT 0.0970 3.1630 0.3450 3.2130 ;
        RECT 0.0970 3.2130 0.1470 3.2160 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.2740 1.4230 0.3340 1.5660 ;
        RECT 0.2210 1.3380 0.3760 1.4230 ;
        RECT 0.0350 1.2880 0.9370 1.3380 ;
        RECT 0.8870 1.3380 0.9370 1.3910 ;
        RECT 0.2740 1.0550 0.3340 1.2880 ;
        RECT 0.7350 1.1200 0.7850 1.2880 ;
        RECT 0.7350 1.3380 0.7850 1.3860 ;
        RECT 0.8870 1.1330 0.9370 1.2880 ;
        RECT 0.8870 1.3910 2.0170 1.4410 ;
    END
  END VDDG

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.5840 1.7020 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.5840 0.0300 ;
        RECT 0.5860 0.0300 0.6360 0.2180 ;
        RECT 0.2790 0.0300 0.3290 0.4410 ;
        RECT 1.5410 0.0300 1.5910 0.3090 ;
        RECT 0.5860 0.2180 0.9370 0.2680 ;
        RECT 1.5410 0.3090 2.0010 0.3590 ;
        RECT 0.7350 0.2680 0.7850 0.4720 ;
        RECT 0.8870 0.2680 0.9370 0.4720 ;
        RECT 1.9510 0.3590 2.0010 0.4830 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 2.5840 3.3740 ;
        RECT 0.4310 3.1430 0.4810 3.3140 ;
        RECT 1.0150 3.0490 1.0650 3.3140 ;
        RECT 1.0150 2.9990 2.1690 3.0490 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 2.6990 2.6650 ;
    LAYER M1 ;
      RECT 0.6950 2.1120 0.8200 2.1620 ;
      RECT 0.6950 2.1620 0.7450 2.5920 ;
      RECT 0.3550 2.5920 0.7450 2.6420 ;
      RECT 0.3550 2.8820 1.6970 2.9320 ;
      RECT 1.3440 2.6040 1.3940 2.8820 ;
      RECT 1.6470 2.6010 1.6970 2.8820 ;
      RECT 1.2510 2.5540 1.3940 2.6040 ;
      RECT 1.6070 2.5510 1.6970 2.6010 ;
      RECT 1.6070 2.3640 1.6570 2.5510 ;
      RECT 1.6070 2.3140 1.7150 2.3640 ;
      RECT 0.3550 2.6420 0.4050 2.8820 ;
      RECT 1.1750 0.3370 1.2650 0.3870 ;
      RECT 1.2150 0.3870 1.2650 1.0100 ;
      RECT 0.4310 1.0100 1.2650 1.0600 ;
      RECT 1.1910 1.0600 1.2410 1.3360 ;
      RECT 0.4310 0.8510 0.4810 1.0100 ;
      RECT 0.4310 0.6010 0.5210 0.6510 ;
      RECT 0.4310 0.4770 0.4810 0.6010 ;
      RECT 0.4310 0.8020 0.5210 0.8510 ;
      RECT 0.4710 0.6510 0.5210 0.8020 ;
      RECT 0.4310 1.0600 0.4810 1.2380 ;
      RECT 1.3430 1.1800 2.2450 1.2300 ;
      RECT 1.3430 1.2300 1.3930 1.3360 ;
      RECT 1.3430 1.0720 1.3930 1.1800 ;
      RECT 1.3150 1.0190 1.3930 1.0720 ;
      RECT 1.3150 0.7680 1.3650 1.0190 ;
      RECT 1.3150 0.7100 1.3930 0.7680 ;
      RECT 1.3430 0.5060 1.3930 0.7100 ;
      RECT 1.3430 0.3770 1.3930 0.4560 ;
      RECT 1.3430 0.4560 1.5610 0.5060 ;
      RECT 1.8100 2.6360 1.9510 2.6860 ;
      RECT 1.8100 2.4640 1.8600 2.6360 ;
      RECT 1.7070 2.4140 1.8600 2.4640 ;
      RECT 1.8100 2.2260 1.8600 2.4140 ;
      RECT 0.9630 2.1760 1.8600 2.2260 ;
      RECT 0.9630 2.2260 1.0130 2.6610 ;
      RECT 0.0350 1.7520 2.1290 1.8080 ;
      RECT 0.6950 1.8080 0.7450 2.0120 ;
      RECT 2.0790 1.8080 2.1290 2.0420 ;
      RECT 0.6950 2.0120 1.4220 2.0620 ;
      RECT 2.0790 2.0420 2.1690 2.0920 ;
      RECT 0.4310 1.8080 0.4810 2.3410 ;
      RECT 1.9510 2.5330 2.3970 2.5830 ;
      RECT 2.2990 2.5830 2.3490 2.8950 ;
      RECT 1.9510 2.0620 2.0010 2.5330 ;
      RECT 1.7800 2.8950 2.3490 2.9450 ;
      RECT 1.7820 2.0120 2.0010 2.0620 ;
      RECT 0.7830 1.5400 2.0930 1.5900 ;
      RECT 1.5550 1.0230 2.3970 1.0730 ;
      RECT 1.1150 3.1010 1.9610 3.1510 ;
      RECT 1.1150 3.1510 1.1650 3.2270 ;
      RECT 1.0390 0.5400 1.1650 0.5900 ;
      RECT 1.0390 0.1680 1.0890 0.5400 ;
      RECT 1.1150 0.5900 1.1650 0.7400 ;
      RECT 1.0390 0.1180 1.4910 0.1680 ;
      RECT 1.0390 0.7400 1.1650 0.7900 ;
      RECT 1.0390 0.7900 1.0890 0.9360 ;
      RECT 1.4710 2.7740 1.5610 2.8240 ;
      RECT 1.4900 2.4100 1.5400 2.7740 ;
      RECT 1.4900 2.3920 1.5450 2.4100 ;
      RECT 1.1510 2.3420 1.5450 2.3920 ;
      RECT 1.1510 2.3920 1.2010 2.7110 ;
      RECT 1.4950 2.3210 1.5450 2.3420 ;
      RECT 0.4910 2.7110 1.2010 2.7610 ;
      RECT 0.5830 0.6400 1.0290 0.6900 ;
      RECT 0.5830 0.6900 0.6330 0.9360 ;
      RECT 0.5830 0.4440 0.6330 0.6400 ;
      RECT 1.4030 3.2010 2.5490 3.2510 ;
      RECT 1.4190 0.8590 1.9410 0.9090 ;
      RECT 1.4190 0.9090 1.4690 0.9460 ;
      RECT 2.0110 2.6800 2.2450 2.7300 ;
      RECT 1.8590 0.5620 2.0930 0.6120 ;
      RECT 0.9470 1.8910 1.1820 1.9410 ;
      RECT 1.4790 1.2860 1.8650 1.3360 ;
    LAYER PO ;
      RECT 1.7330 1.7550 1.7630 2.4920 ;
      RECT 0.6690 1.7550 0.6990 3.2820 ;
      RECT 1.7330 2.6520 1.7630 3.2820 ;
      RECT 0.3650 1.7400 0.3950 3.2820 ;
      RECT 1.2770 0.0900 1.3070 0.5640 ;
      RECT 0.8210 1.7550 0.8510 3.2820 ;
      RECT 1.8850 0.7800 1.9150 3.2820 ;
      RECT 0.5170 0.0900 0.5470 1.6280 ;
      RECT 1.5810 0.0900 1.6110 1.6280 ;
      RECT 0.9730 0.0900 1.0030 1.6280 ;
      RECT 1.4290 0.0900 1.4590 1.6280 ;
      RECT 0.8210 0.0900 0.8510 1.6280 ;
      RECT 1.7330 0.0900 1.7630 1.6280 ;
      RECT 0.6690 0.0900 0.6990 1.6280 ;
      RECT 2.0370 0.0900 2.0670 1.6280 ;
      RECT 1.1250 0.0900 1.1550 3.2820 ;
      RECT 0.3650 0.0900 0.3950 1.6280 ;
      RECT 1.5810 1.7550 1.6110 3.2820 ;
      RECT 1.4290 1.7550 1.4590 3.2820 ;
      RECT 0.5170 1.7400 0.5470 3.2820 ;
      RECT 2.0370 1.7550 2.0670 3.2820 ;
      RECT 2.4930 0.0900 2.5230 3.2820 ;
      RECT 1.8850 0.0900 1.9150 0.6400 ;
      RECT 1.2770 1.7550 1.3070 3.2820 ;
      RECT 0.2130 0.2490 0.2430 3.2820 ;
      RECT 2.1890 0.0900 2.2190 3.2820 ;
      RECT 0.9730 2.5610 1.0030 3.2820 ;
      RECT 0.0610 0.2490 0.0910 3.2820 ;
      RECT 2.3410 0.0900 2.3710 3.2820 ;
      RECT 0.9730 1.7550 1.0030 2.3580 ;
      RECT 1.2770 1.0120 1.3070 1.6280 ;
  END
END AODFFNARX1_LVT

MACRO AODFFNARX2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.888 BY 3.344 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8570 1.4630 1.0290 1.5920 ;
    END
    ANTENNAGATEAREA 0.0342 ;
  END CLK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 0.6970 0.6630 0.7020 ;
        RECT 0.5530 0.7020 0.7250 0.7520 ;
        RECT 0.5530 0.7520 0.6630 0.8140 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END D

  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.0270 0.1080 2.8530 0.1580 ;
        RECT 2.0270 0.0970 2.1830 0.1080 ;
        RECT 2.0270 0.1580 2.1830 0.2070 ;
    END
    ANTENNAGATEAREA 0.0441 ;
  END RSTB

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0970 3.1430 0.2070 3.2530 ;
        RECT 0.1150 3.0800 0.1650 3.1430 ;
        RECT 0.1150 3.0300 0.4810 3.0800 ;
        RECT 0.1150 2.4320 0.1650 3.0300 ;
        RECT 0.4310 3.0800 0.4810 3.2020 ;
        RECT 0.1150 2.3820 0.4810 2.4320 ;
        RECT 0.4310 1.8780 0.4810 2.3820 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2390 2.4960 0.7850 2.5460 ;
        RECT 0.7350 1.8880 0.7850 2.4960 ;
        RECT 0.2390 2.5460 0.2890 2.8390 ;
        RECT 0.2390 2.8390 0.3590 2.9200 ;
        RECT 0.2390 2.9200 0.7850 2.9700 ;
        RECT 0.7350 2.9700 0.7850 3.2020 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q

  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.5780 1.4230 0.6380 1.5660 ;
        RECT 0.5250 1.3380 0.6800 1.4230 ;
        RECT 0.0350 1.2880 1.2410 1.3380 ;
        RECT 1.1910 1.3380 1.2410 1.3910 ;
        RECT 0.5780 1.0550 0.6380 1.2880 ;
        RECT 1.0390 1.3380 1.0890 1.3860 ;
        RECT 1.0390 1.1200 1.0890 1.2880 ;
        RECT 1.1910 1.1330 1.2410 1.2880 ;
        RECT 1.1910 1.3910 2.3210 1.4410 ;
    END
  END VDDG

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.8880 1.7020 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.8880 0.0300 ;
        RECT 0.8900 0.0300 0.9400 0.2180 ;
        RECT 0.5830 0.0300 0.6330 0.4410 ;
        RECT 1.8450 0.0300 1.8950 0.3090 ;
        RECT 0.8900 0.2180 1.2410 0.2680 ;
        RECT 1.8450 0.3090 2.3050 0.3590 ;
        RECT 1.0390 0.2680 1.0890 0.4720 ;
        RECT 1.1910 0.2680 1.2410 0.4720 ;
        RECT 2.2550 0.3590 2.3050 0.4830 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 3.3140 2.8880 3.3740 ;
        RECT 0.5830 3.0380 0.6330 3.3140 ;
        RECT 0.2790 3.1300 0.3290 3.3140 ;
        RECT 0.8870 2.9270 0.9370 3.3140 ;
        RECT 1.3190 3.0490 1.3690 3.3140 ;
        RECT 1.3190 2.9990 2.4730 3.0490 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 3.0030 2.6650 ;
    LAYER M1 ;
      RECT 1.6480 2.8820 2.0010 2.9320 ;
      RECT 1.6480 2.8460 1.6980 2.8820 ;
      RECT 1.9510 2.6010 2.0010 2.8820 ;
      RECT 0.5260 2.7960 1.6980 2.8460 ;
      RECT 1.9110 2.5510 2.0010 2.6010 ;
      RECT 1.6480 2.6040 1.6980 2.7960 ;
      RECT 1.9110 2.3640 1.9610 2.5510 ;
      RECT 1.5550 2.5540 1.6980 2.6040 ;
      RECT 1.9110 2.3140 2.0190 2.3640 ;
      RECT 0.9990 2.1620 1.0490 2.5960 ;
      RECT 0.9990 2.1120 1.1240 2.1620 ;
      RECT 0.5260 2.5960 1.0490 2.6460 ;
      RECT 0.5260 2.8460 0.5760 2.8470 ;
      RECT 0.5260 2.7460 0.5760 2.7960 ;
      RECT 0.3390 2.6960 0.5760 2.7460 ;
      RECT 0.5260 2.6460 0.5760 2.6960 ;
      RECT 1.4790 0.3370 1.5690 0.3870 ;
      RECT 1.5190 0.3870 1.5690 1.0100 ;
      RECT 0.7350 1.0100 1.5690 1.0600 ;
      RECT 1.4950 1.0600 1.5450 1.3360 ;
      RECT 0.7350 0.8510 0.7850 1.0100 ;
      RECT 0.7350 0.6010 0.8250 0.6510 ;
      RECT 0.7350 0.4770 0.7850 0.6010 ;
      RECT 0.7350 0.8020 0.8250 0.8510 ;
      RECT 0.7750 0.6510 0.8250 0.8020 ;
      RECT 0.7350 1.0600 0.7850 1.2380 ;
      RECT 1.6470 1.1800 2.5490 1.2300 ;
      RECT 1.6470 1.2300 1.6970 1.3360 ;
      RECT 1.6470 1.0720 1.6970 1.1800 ;
      RECT 1.6190 1.0190 1.6970 1.0720 ;
      RECT 1.6190 0.7680 1.6690 1.0190 ;
      RECT 1.6190 0.7100 1.6970 0.7680 ;
      RECT 1.6470 0.5060 1.6970 0.7100 ;
      RECT 1.6470 0.3770 1.6970 0.4560 ;
      RECT 1.6470 0.4560 1.8650 0.5060 ;
      RECT 1.2510 1.8910 1.4860 1.9410 ;
      RECT 1.4190 3.1040 2.2650 3.1540 ;
      RECT 1.4190 3.1540 1.4690 3.2270 ;
      RECT 1.3430 0.5400 1.4690 0.5900 ;
      RECT 1.3430 0.1680 1.3930 0.5400 ;
      RECT 1.4190 0.5900 1.4690 0.7400 ;
      RECT 1.3430 0.1180 1.7950 0.1680 ;
      RECT 1.3430 0.7400 1.4690 0.7900 ;
      RECT 1.3430 0.7900 1.3930 0.9360 ;
      RECT 2.3830 2.0420 2.4730 2.0920 ;
      RECT 2.3830 1.8080 2.4330 2.0420 ;
      RECT 0.0350 1.7520 2.4330 1.8080 ;
      RECT 0.8870 1.8080 0.9370 2.4380 ;
      RECT 0.9990 1.8080 1.0490 2.0120 ;
      RECT 0.9990 2.0120 1.7260 2.0620 ;
      RECT 0.5830 1.8080 0.6330 2.3900 ;
      RECT 0.2790 1.8080 0.3290 2.2980 ;
      RECT 2.0860 2.0120 2.3050 2.0620 ;
      RECT 2.2550 2.0620 2.3050 2.5330 ;
      RECT 2.2550 2.5330 2.7010 2.5830 ;
      RECT 2.6030 2.5830 2.6530 2.8950 ;
      RECT 2.0840 2.8950 2.6530 2.9450 ;
      RECT 1.7830 1.2860 2.1690 1.3360 ;
      RECT 2.1140 2.6360 2.2550 2.6860 ;
      RECT 2.1140 2.4640 2.1640 2.6360 ;
      RECT 2.0110 2.4140 2.1640 2.4640 ;
      RECT 2.1140 2.2260 2.1640 2.4140 ;
      RECT 1.2670 2.1760 2.1640 2.2260 ;
      RECT 1.2670 2.2260 1.3170 2.6460 ;
      RECT 1.0990 1.5400 2.3970 1.5900 ;
      RECT 1.8590 1.0230 2.7010 1.0730 ;
      RECT 1.7750 2.7740 1.8650 2.8240 ;
      RECT 1.7940 2.4100 1.8440 2.7740 ;
      RECT 1.7940 2.3920 1.8490 2.4100 ;
      RECT 1.4550 2.3420 1.8490 2.3920 ;
      RECT 1.4550 2.3920 1.5050 2.6960 ;
      RECT 1.7990 2.3210 1.8490 2.3420 ;
      RECT 0.6430 2.6960 1.5050 2.7460 ;
      RECT 0.8870 0.6400 1.3330 0.6900 ;
      RECT 0.8870 0.6900 0.9370 0.9360 ;
      RECT 0.8870 0.4440 0.9370 0.6400 ;
      RECT 1.7070 3.2040 2.8530 3.2540 ;
      RECT 1.7230 0.8590 2.2450 0.9090 ;
      RECT 1.7230 0.9090 1.7730 0.9460 ;
      RECT 2.3150 2.6800 2.5490 2.7300 ;
      RECT 2.1630 0.5620 2.3970 0.6120 ;
    LAYER PO ;
      RECT 0.9730 1.7400 1.0030 3.2820 ;
      RECT 0.8210 1.7400 0.8510 3.2820 ;
      RECT 0.6690 1.7400 0.6990 3.2820 ;
      RECT 0.5170 0.2490 0.5470 3.2820 ;
      RECT 0.0610 0.0900 0.0910 3.2820 ;
      RECT 0.3650 1.7400 0.3950 3.2820 ;
      RECT 0.2130 1.7400 0.2430 3.2820 ;
      RECT 0.2130 0.0900 0.2430 1.6280 ;
      RECT 2.1890 0.0900 2.2190 0.6400 ;
      RECT 1.5810 1.7550 1.6110 3.2820 ;
      RECT 2.4930 0.0900 2.5230 3.2820 ;
      RECT 1.2770 2.5460 1.3070 3.2820 ;
      RECT 2.6450 0.0900 2.6750 3.2820 ;
      RECT 1.2770 1.7550 1.3070 2.3580 ;
      RECT 1.5810 1.0120 1.6110 1.6280 ;
      RECT 2.0370 1.7550 2.0670 2.4920 ;
      RECT 2.0370 2.6520 2.0670 3.2820 ;
      RECT 1.5810 0.0900 1.6110 0.5640 ;
      RECT 1.1250 1.7550 1.1550 3.2820 ;
      RECT 2.1890 0.7800 2.2190 3.2820 ;
      RECT 0.8210 0.0900 0.8510 1.6280 ;
      RECT 1.8850 0.0900 1.9150 1.6280 ;
      RECT 1.2770 0.0900 1.3070 1.6280 ;
      RECT 1.7330 0.0900 1.7630 1.6280 ;
      RECT 1.1250 0.0900 1.1550 1.6280 ;
      RECT 2.0370 0.0900 2.0670 1.6280 ;
      RECT 0.9730 0.0900 1.0030 1.6280 ;
      RECT 2.3410 0.0900 2.3710 1.6280 ;
      RECT 1.4290 0.0900 1.4590 3.2820 ;
      RECT 0.6690 0.0900 0.6990 1.6280 ;
      RECT 1.8850 1.7550 1.9150 3.2820 ;
      RECT 0.3650 0.2490 0.3950 1.6210 ;
      RECT 1.7330 1.7550 1.7630 3.2820 ;
      RECT 2.3410 1.7550 2.3710 3.2820 ;
      RECT 2.7970 0.0900 2.8270 3.2820 ;
  END
END AODFFNARX2_LVT

MACRO AOI21X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.824 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.8240 0.0300 ;
        RECT 1.0390 0.0300 1.0890 0.5620 ;
        RECT 1.3430 0.0300 1.3930 0.4890 ;
        RECT 0.2790 0.0300 0.3290 0.2880 ;
        RECT 0.2790 0.2880 0.7850 0.3380 ;
        RECT 0.7350 0.3380 0.7850 0.5620 ;
        RECT 0.2790 0.3380 0.3290 0.5620 ;
    END
  END VSS

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4650 1.1610 1.5750 1.2710 ;
        RECT 1.4950 1.2710 1.5450 1.5540 ;
        RECT 1.4950 0.8530 1.5450 1.1610 ;
        RECT 1.4950 0.8030 1.5850 0.8530 ;
        RECT 1.5350 0.5010 1.5850 0.8030 ;
        RECT 1.4950 0.4300 1.5850 0.5010 ;
        RECT 1.4950 0.1140 1.5450 0.4300 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7050 0.4210 0.8150 ;
    END
    ANTENNAGATEAREA 0.0243 ;
  END A2

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.8240 1.7020 ;
        RECT 0.5830 1.1720 0.6330 1.6420 ;
        RECT 0.2790 1.0280 0.3290 1.6420 ;
        RECT 1.0390 1.0000 1.0890 1.6420 ;
        RECT 1.3420 1.1040 1.3920 1.6420 ;
    END
  END VDD

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 0.0970 0.8770 0.2070 ;
    END
    ANTENNAGATEAREA 0.0228 ;
  END A3

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4920 0.8570 0.6630 0.9670 ;
    END
    ANTENNAGATEAREA 0.0243 ;
  END A1
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.9390 1.7870 ;
    LAYER M1 ;
      RECT 0.5830 0.3880 0.6330 0.7570 ;
      RECT 0.8870 0.8070 0.9370 1.5630 ;
      RECT 0.8870 0.3880 0.9370 0.7570 ;
      RECT 0.5830 0.7570 1.1810 0.8070 ;
      RECT 1.1910 0.6230 1.4850 0.6730 ;
      RECT 1.3460 0.6730 1.3960 0.9610 ;
      RECT 1.1910 0.9610 1.3960 1.0110 ;
      RECT 1.1910 0.3880 1.2410 0.6230 ;
      RECT 1.1910 1.0110 1.2410 1.5230 ;
      RECT 0.7350 1.0770 0.7850 1.5200 ;
      RECT 0.4310 1.0270 0.7850 1.0770 ;
      RECT 0.4310 1.0770 0.4810 1.5250 ;
    LAYER PO ;
      RECT 1.5810 0.0630 1.6110 1.6040 ;
      RECT 0.2130 0.0640 0.2430 1.6130 ;
      RECT 1.4290 0.0640 1.4590 1.6040 ;
      RECT 0.9730 0.0640 1.0030 1.6130 ;
      RECT 1.2770 0.0590 1.3070 1.6130 ;
      RECT 0.5170 0.0640 0.5470 1.6130 ;
      RECT 0.0610 0.0640 0.0910 1.6130 ;
      RECT 1.7330 0.0630 1.7630 1.6040 ;
      RECT 0.3650 0.0590 0.3950 1.6130 ;
      RECT 0.8210 0.0590 0.8510 1.6130 ;
      RECT 0.6690 0.0640 0.6990 1.6130 ;
      RECT 1.1250 0.0590 1.1550 1.6130 ;
  END
END AOI21X1_LVT

MACRO AND2X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.216 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8870 0.1170 0.9370 0.5520 ;
        RECT 0.8870 0.5520 1.0450 0.5530 ;
        RECT 0.8870 0.5530 1.1190 0.6020 ;
        RECT 0.9740 0.6020 1.1190 0.6630 ;
        RECT 0.9740 0.6630 1.0240 0.8590 ;
        RECT 0.8870 0.8590 1.0240 0.9090 ;
        RECT 0.8870 0.9090 0.9370 1.5590 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 0.8870 0.5730 0.9370 ;
        RECT 0.4010 0.8570 0.5110 0.8870 ;
        RECT 0.4010 0.9370 0.5110 0.9670 ;
    END
    ANTENNAGATEAREA 0.0243 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7350 0.4210 0.7850 ;
        RECT 0.2490 0.7050 0.3590 0.7350 ;
        RECT 0.2490 0.7850 0.3590 0.8150 ;
    END
    ANTENNAGATEAREA 0.0243 ;
  END A2

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.2160 1.7020 ;
        RECT 0.7350 0.8930 0.7850 1.6420 ;
        RECT 0.4310 1.3630 0.4810 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.2160 0.0300 ;
        RECT 0.7350 0.0300 0.7850 0.5030 ;
        RECT 0.2790 0.0300 0.3290 0.4790 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.3310 1.7730 ;
    LAYER M1 ;
      RECT 0.5830 0.6560 0.8770 0.7060 ;
      RECT 0.2790 1.0940 0.3290 1.5690 ;
      RECT 0.6240 0.6560 0.6740 1.1430 ;
      RECT 0.5830 0.1060 0.6330 0.6960 ;
      RECT 0.3040 1.0940 0.6720 1.1440 ;
      RECT 0.5830 1.1190 0.6330 1.5690 ;
    LAYER PO ;
      RECT 0.3650 0.0710 0.3950 1.6040 ;
      RECT 0.5170 0.0710 0.5470 1.6040 ;
      RECT 0.2130 0.0710 0.2430 1.6040 ;
      RECT 0.0610 0.0710 0.0910 1.6040 ;
      RECT 0.9730 0.0720 1.0030 1.6040 ;
      RECT 1.1250 0.0720 1.1550 1.6040 ;
      RECT 0.8210 0.0720 0.8510 1.6060 ;
      RECT 0.6690 0.0710 0.6990 1.6040 ;
  END
END AND2X1_LVT

MACRO AND2X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.368 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1310 0.5530 1.2710 0.6630 ;
        RECT 0.7350 0.5030 1.1810 0.5530 ;
        RECT 1.1310 0.6630 1.1810 0.7030 ;
        RECT 0.7350 0.1300 0.7850 0.5030 ;
        RECT 1.0390 0.1300 1.0890 0.5030 ;
        RECT 0.7350 0.7030 1.1810 0.7530 ;
        RECT 1.0390 0.7530 1.0890 1.5440 ;
        RECT 0.7350 0.7530 0.7850 1.5440 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4910 0.7350 0.6630 0.7850 ;
        RECT 0.5530 0.7050 0.6630 0.7350 ;
        RECT 0.5530 0.7850 0.6630 0.8150 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7050 0.3590 0.7350 ;
        RECT 0.2490 0.7350 0.4210 0.7850 ;
        RECT 0.2490 0.7850 0.3590 0.8150 ;
    END
    ANTENNAGATEAREA 0.024 ;
  END A2

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.3680 1.7020 ;
        RECT 0.8870 0.8180 0.9370 1.6420 ;
        RECT 0.4310 1.1950 0.4810 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.3680 0.0300 ;
        RECT 0.8870 0.0300 0.9370 0.3980 ;
        RECT 0.2790 0.0300 0.3290 0.4790 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.4830 1.7730 ;
    LAYER M1 ;
      RECT 0.1490 0.6030 1.0290 0.6530 ;
      RECT 0.1490 0.6080 0.1990 0.9150 ;
      RECT 0.2790 0.8650 0.3290 1.5530 ;
      RECT 0.5830 0.1210 0.6330 0.6470 ;
      RECT 0.5830 0.8890 0.6330 1.5530 ;
      RECT 0.1500 0.8650 0.6330 0.9150 ;
    LAYER PO ;
      RECT 0.9730 0.0720 1.0030 1.6040 ;
      RECT 1.1250 0.0720 1.1550 1.6030 ;
      RECT 0.8210 0.0720 0.8510 1.6040 ;
      RECT 0.6690 0.0710 0.6990 1.6030 ;
      RECT 0.3650 0.0710 0.3950 1.6030 ;
      RECT 0.5170 0.0710 0.5470 1.6030 ;
      RECT 0.2130 0.0710 0.2430 1.6030 ;
      RECT 0.0610 0.0710 0.0910 1.6030 ;
      RECT 1.2770 0.0720 1.3070 1.6100 ;
  END
END AND2X2_LVT

MACRO AND2X4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.672 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7370 0.4210 0.7870 ;
        RECT 0.2490 0.7060 0.3590 0.7370 ;
        RECT 0.2490 0.7870 0.3590 0.8160 ;
    END
    ANTENNAGATEAREA 0.0234 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4910 0.7370 0.6630 0.7870 ;
        RECT 0.5530 0.7870 0.6630 0.8170 ;
        RECT 0.5530 0.7070 0.6630 0.7370 ;
    END
    ANTENNAGATEAREA 0.0234 ;
  END A1

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.6720 0.0300 ;
        RECT 1.1910 0.0300 1.2410 0.3980 ;
        RECT 0.2790 0.0300 0.3290 0.4800 ;
        RECT 0.8870 0.0300 0.9370 0.3980 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.6720 1.7020 ;
        RECT 0.4310 1.1960 0.4810 1.6420 ;
        RECT 1.1910 0.8180 1.2410 1.6420 ;
        RECT 0.8870 0.8180 0.9370 1.6420 ;
    END
  END VDD

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4280 0.5330 1.4780 0.5530 ;
        RECT 1.4280 0.5530 1.5750 0.6630 ;
        RECT 0.7350 0.4830 1.4780 0.5330 ;
        RECT 1.4280 0.6630 1.4780 0.7090 ;
        RECT 1.3430 0.1320 1.3930 0.4830 ;
        RECT 1.0390 0.1300 1.0890 0.4830 ;
        RECT 0.7350 0.1300 0.7850 0.4830 ;
        RECT 0.7350 0.7090 1.4780 0.7590 ;
        RECT 1.3430 0.7590 1.3930 1.5440 ;
        RECT 1.0390 0.7590 1.0890 1.5440 ;
        RECT 0.7350 0.7590 0.7850 1.5440 ;
    END
    ANTENNADIFFAREA 0.3972 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.7870 1.7730 ;
    LAYER M1 ;
      RECT 0.1490 0.5910 1.3330 0.6410 ;
      RECT 0.1490 0.6170 0.1990 0.9170 ;
      RECT 0.2790 0.8670 0.3290 1.5540 ;
      RECT 0.5830 0.1220 0.6330 0.6410 ;
      RECT 0.5830 0.8920 0.6330 1.5540 ;
      RECT 0.1490 0.8670 0.6330 0.9170 ;
    LAYER PO ;
      RECT 0.2130 0.0710 0.2430 1.6040 ;
      RECT 0.5170 0.0710 0.5470 1.6040 ;
      RECT 0.3650 0.0710 0.3950 1.6040 ;
      RECT 0.6690 0.0710 0.6990 1.6040 ;
      RECT 0.8210 0.0720 0.8510 1.6040 ;
      RECT 1.4290 0.0720 1.4590 1.6040 ;
      RECT 1.5810 0.0720 1.6110 1.6040 ;
      RECT 1.2770 0.0720 1.3070 1.6040 ;
      RECT 1.1250 0.0720 1.1550 1.6040 ;
      RECT 0.9730 0.0720 1.0030 1.6040 ;
      RECT 0.0610 0.0710 0.0910 1.6040 ;
  END
END AND2X4_LVT

MACRO AND3X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.368 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 0.7370 0.7250 0.7870 ;
        RECT 0.5530 0.7070 0.6630 0.7370 ;
        RECT 0.5530 0.7870 0.6630 0.8170 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0390 0.4800 1.1660 0.5300 ;
        RECT 1.0390 0.1210 1.0890 0.4800 ;
        RECT 1.1160 0.5300 1.1660 0.7050 ;
        RECT 1.1160 0.7050 1.2710 0.7650 ;
        RECT 1.0390 0.7650 1.2710 0.8150 ;
        RECT 1.0390 0.8150 1.0890 1.5440 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 1.0410 0.5730 1.0910 ;
        RECT 0.4010 1.0110 0.5110 1.0410 ;
        RECT 0.4010 1.0910 0.5110 1.1210 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END A2

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.3680 0.0300 ;
        RECT 0.2790 0.0300 0.3290 0.4790 ;
        RECT 0.8870 0.0300 0.9370 0.4790 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.3680 1.7020 ;
        RECT 0.8870 0.8180 0.9370 1.6420 ;
        RECT 0.2790 1.2850 0.3290 1.6420 ;
        RECT 0.5830 1.2850 0.6330 1.6420 ;
    END
  END VDD

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7070 0.3590 0.7370 ;
        RECT 0.2490 0.7370 0.4210 0.7870 ;
        RECT 0.2490 0.7870 0.3590 0.8170 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END A3
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.4830 1.7730 ;
    LAYER M1 ;
      RECT 0.7840 0.6580 1.0480 0.7080 ;
      RECT 0.4310 1.1840 0.4810 1.5530 ;
      RECT 0.7350 0.1210 0.7850 0.6140 ;
      RECT 0.4560 1.1840 0.8090 1.2340 ;
      RECT 0.7350 1.1870 0.7850 1.5530 ;
      RECT 0.7350 0.5650 0.8080 0.6150 ;
      RECT 0.7750 0.5650 0.8250 1.2340 ;
    LAYER PO ;
      RECT 1.1250 0.0720 1.1550 1.6030 ;
      RECT 1.2770 0.0720 1.3070 1.6030 ;
      RECT 0.9730 0.0710 1.0030 1.6040 ;
      RECT 0.0610 0.0710 0.0910 1.6030 ;
      RECT 0.8210 0.0710 0.8510 1.6030 ;
      RECT 0.2130 0.0710 0.2430 1.6030 ;
      RECT 0.5170 0.0710 0.5470 1.6030 ;
      RECT 0.3650 0.0710 0.3950 1.6030 ;
      RECT 0.6690 0.0710 0.6990 1.6030 ;
  END
END AND3X1_LVT

MACRO AND3X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.52 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2780 0.5530 1.4230 0.6630 ;
        RECT 1.2780 0.5290 1.3280 0.5530 ;
        RECT 1.2780 0.6630 1.3280 0.7140 ;
        RECT 0.8870 0.4790 1.3280 0.5290 ;
        RECT 0.8870 0.7140 1.3280 0.7640 ;
        RECT 0.8870 0.1290 0.9370 0.4790 ;
        RECT 1.1910 0.1290 1.2410 0.4790 ;
        RECT 1.1910 0.7640 1.2410 1.5440 ;
        RECT 0.8870 0.7640 0.9370 1.5440 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END Y

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7350 0.4210 0.7850 ;
        RECT 0.2490 0.7050 0.3590 0.7350 ;
        RECT 0.2490 0.7850 0.3590 0.8150 ;
    END
    ANTENNAGATEAREA 0.0198 ;
  END A3

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.5200 1.7020 ;
        RECT 1.0390 0.8140 1.0890 1.6420 ;
        RECT 0.5830 1.3790 0.6330 1.6420 ;
        RECT 0.2790 1.3790 0.3290 1.6420 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.5200 0.0300 ;
        RECT 1.0410 0.0300 1.0910 0.3980 ;
        RECT 0.2790 0.0300 0.3290 0.4790 ;
    END
  END VSS

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 1.0090 0.5110 1.0390 ;
        RECT 0.4010 1.0390 0.5730 1.0890 ;
        RECT 0.4010 1.0890 0.5110 1.1190 ;
    END
    ANTENNAGATEAREA 0.0198 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 0.7050 0.6630 0.7350 ;
        RECT 0.5530 0.7350 0.7250 0.7850 ;
        RECT 0.5530 0.7850 0.6630 0.8150 ;
    END
    ANTENNAGATEAREA 0.0198 ;
  END A1
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.6350 1.7730 ;
    LAYER M1 ;
      RECT 0.7350 0.6140 1.1810 0.6640 ;
      RECT 0.7350 0.1210 0.7850 0.6420 ;
      RECT 0.7350 1.1870 0.7850 1.5530 ;
      RECT 0.4560 1.1870 0.8250 1.2370 ;
      RECT 0.7750 0.6140 0.8250 1.2110 ;
      RECT 0.4310 1.1870 0.4810 1.5530 ;
    LAYER PO ;
      RECT 1.1250 0.0710 1.1550 1.6040 ;
      RECT 1.2770 0.0720 1.3070 1.6030 ;
      RECT 0.9730 0.0710 1.0030 1.6040 ;
      RECT 1.4290 0.0720 1.4590 1.6030 ;
      RECT 0.6690 0.0710 0.6990 1.6030 ;
      RECT 0.3650 0.0710 0.3950 1.6030 ;
      RECT 0.5170 0.0710 0.5470 1.6030 ;
      RECT 0.2130 0.0710 0.2430 1.6030 ;
      RECT 0.8210 0.0710 0.8510 1.6030 ;
      RECT 0.0610 0.0710 0.0910 1.6030 ;
  END
END AND3X2_LVT

MACRO AND3X4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.824 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4950 0.1150 1.5450 0.5220 ;
        RECT 0.8870 0.5220 1.6660 0.5530 ;
        RECT 1.1910 0.1150 1.2410 0.5220 ;
        RECT 0.8870 0.1150 0.9370 0.5220 ;
        RECT 0.8870 0.5530 1.7360 0.5720 ;
        RECT 1.6160 0.5720 1.7360 0.6630 ;
        RECT 1.6160 0.6630 1.6660 0.7220 ;
        RECT 0.8870 0.7220 1.6660 0.7720 ;
        RECT 1.4950 0.7720 1.5450 1.5590 ;
        RECT 1.1910 0.7720 1.2410 1.5590 ;
        RECT 0.8870 0.7720 0.9370 1.5590 ;
    END
    ANTENNADIFFAREA 0.3972 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 0.7350 0.7250 0.7850 ;
        RECT 0.5530 0.7050 0.6630 0.7350 ;
        RECT 0.5530 0.7850 0.6630 0.8150 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 1.0090 0.5110 1.0390 ;
        RECT 0.4010 1.0390 0.5730 1.0890 ;
        RECT 0.4010 1.0890 0.5110 1.1190 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END A2

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.8240 0.0300 ;
        RECT 1.3430 0.0300 1.3930 0.4130 ;
        RECT 1.0390 0.0300 1.0890 0.4130 ;
        RECT 0.2790 0.0300 0.3290 0.4790 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.8240 1.7020 ;
        RECT 1.3430 0.9100 1.3930 1.6420 ;
        RECT 1.0390 0.9100 1.0890 1.6420 ;
        RECT 0.2790 1.3790 0.3290 1.6420 ;
        RECT 0.5830 1.3790 0.6330 1.6420 ;
    END
  END VDD

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7350 0.4210 0.7850 ;
        RECT 0.2490 0.7050 0.3590 0.7350 ;
        RECT 0.2490 0.7850 0.3590 0.8150 ;
    END
    ANTENNAGATEAREA 0.0204 ;
  END A3
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.9390 1.7730 ;
    LAYER M1 ;
      RECT 0.7840 0.6220 1.4850 0.6720 ;
      RECT 0.4310 1.1850 0.4810 1.5530 ;
      RECT 0.7800 0.5710 0.8300 1.2100 ;
      RECT 0.7350 0.1210 0.7850 0.6140 ;
      RECT 0.4560 1.1850 0.8300 1.2350 ;
      RECT 0.7350 1.1850 0.7850 1.5530 ;
      RECT 0.7350 0.5690 0.8300 0.6190 ;
    LAYER PO ;
      RECT 0.9730 0.0720 1.0030 1.6040 ;
      RECT 1.5810 0.0720 1.6110 1.6030 ;
      RECT 1.7330 0.0720 1.7630 1.6030 ;
      RECT 1.4290 0.0720 1.4590 1.6040 ;
      RECT 1.2770 0.0720 1.3070 1.6040 ;
      RECT 1.1250 0.0720 1.1550 1.6040 ;
      RECT 0.0610 0.0710 0.0910 1.6030 ;
      RECT 0.8210 0.0710 0.8510 1.6030 ;
      RECT 0.2130 0.0710 0.2430 1.6030 ;
      RECT 0.5170 0.0710 0.5470 1.6030 ;
      RECT 0.3650 0.0710 0.3950 1.6030 ;
      RECT 0.6690 0.0710 0.6990 1.6030 ;
  END
END AND3X4_LVT

MACRO AND4X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.52 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1910 0.1170 1.2410 0.5510 ;
        RECT 1.1910 0.5510 1.3150 0.5530 ;
        RECT 1.1910 0.5530 1.4330 0.6010 ;
        RECT 1.2900 0.6010 1.4330 0.6630 ;
        RECT 1.2900 0.6630 1.3400 0.7550 ;
        RECT 1.1910 0.7550 1.3400 0.8050 ;
        RECT 1.1910 0.8050 1.2410 1.5570 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 1.0390 0.8770 1.0890 ;
        RECT 0.7050 1.0090 0.8150 1.0390 ;
        RECT 0.7050 1.0890 0.8150 1.1190 ;
    END
    ANTENNAGATEAREA 0.0183 ;
  END A1

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 1.0390 0.5730 1.0890 ;
        RECT 0.4010 1.0090 0.5110 1.0390 ;
        RECT 0.4010 1.0890 0.5110 1.1190 ;
    END
    ANTENNAGATEAREA 0.0183 ;
  END A3

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7050 0.3590 0.7350 ;
        RECT 0.2490 0.7350 0.4210 0.7850 ;
        RECT 0.2490 0.7850 0.3590 0.8150 ;
    END
    ANTENNAGATEAREA 0.0183 ;
  END A4

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.5200 0.0300 ;
        RECT 1.0390 0.0300 1.0890 0.4880 ;
        RECT 0.2790 0.0300 0.3290 0.4790 ;
    END
  END VSS

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 0.7050 0.6630 0.7350 ;
        RECT 0.5530 0.7350 0.7250 0.7850 ;
        RECT 0.5530 0.7850 0.6630 0.8150 ;
    END
    ANTENNAGATEAREA 0.0183 ;
  END A2

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.5200 1.7020 ;
        RECT 1.0390 0.8310 1.0890 1.6420 ;
        RECT 0.7350 1.3820 0.7850 1.6420 ;
        RECT 0.4310 1.3820 0.4810 1.6420 ;
    END
  END VDD
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.6350 1.7730 ;
    LAYER M1 ;
      RECT 0.9700 0.6510 1.1810 0.7000 ;
      RECT 0.9700 0.6500 1.1410 0.6510 ;
      RECT 0.2790 1.2600 0.3290 1.5560 ;
      RECT 0.5830 1.2860 0.6330 1.5560 ;
      RECT 0.8870 0.6220 0.9700 0.6720 ;
      RECT 0.8870 0.1210 0.9370 0.6470 ;
      RECT 0.2790 1.2630 0.9770 1.3130 ;
      RECT 0.8870 1.2760 0.9370 1.5560 ;
      RECT 0.9270 0.6220 0.9770 1.2880 ;
    LAYER PO ;
      RECT 1.2770 0.0720 1.3070 1.6090 ;
      RECT 1.4290 0.0720 1.4590 1.6090 ;
      RECT 1.1250 0.0720 1.1550 1.6090 ;
      RECT 0.9730 0.0710 1.0030 1.6090 ;
      RECT 0.6690 0.0710 0.6990 1.6090 ;
      RECT 0.3650 0.0710 0.3950 1.6090 ;
      RECT 0.5170 0.0710 0.5470 1.6090 ;
      RECT 0.2130 0.0710 0.2430 1.6090 ;
      RECT 0.8210 0.0710 0.8510 1.6090 ;
      RECT 0.0610 0.0710 0.0910 1.6090 ;
  END
END AND4X1_LVT

MACRO AND4X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.28 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 0.7350 0.7250 0.7850 ;
        RECT 0.5530 0.7050 0.6630 0.7350 ;
        RECT 0.5530 0.7850 0.6630 0.8150 ;
    END
    ANTENNAGATEAREA 0.0165 ;
  END A2

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.2800 0.0300 ;
        RECT 1.6470 0.0300 1.6970 0.4860 ;
        RECT 1.3430 0.0300 1.3930 0.3020 ;
        RECT 1.9510 0.0300 2.0010 0.4860 ;
        RECT 1.0390 0.0300 1.0890 0.3040 ;
        RECT 0.2790 0.0300 0.3290 0.4790 ;
    END
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.2800 1.7020 ;
        RECT 1.6470 0.8230 1.6970 1.6420 ;
        RECT 1.9510 0.9150 2.0010 1.6420 ;
        RECT 1.3430 1.0990 1.3930 1.6420 ;
        RECT 0.7350 1.3820 0.7850 1.6420 ;
        RECT 1.0390 1.1990 1.0890 1.6420 ;
        RECT 0.4310 1.3780 0.4810 1.6420 ;
    END
  END VDD

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7050 0.3590 0.7350 ;
        RECT 0.2490 0.7350 0.4210 0.7850 ;
        RECT 0.2490 0.7850 0.3590 0.8150 ;
    END
    ANTENNAGATEAREA 0.0165 ;
  END A4

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 1.0090 0.5110 1.0390 ;
        RECT 0.4010 1.0390 0.5730 1.0890 ;
        RECT 0.4010 1.0890 0.5110 1.1190 ;
    END
    ANTENNAGATEAREA 0.0165 ;
  END A3

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 1.0090 0.8150 1.0390 ;
        RECT 0.7050 1.0390 0.8770 1.0890 ;
        RECT 0.7050 1.0890 0.8150 1.1190 ;
    END
    ANTENNAGATEAREA 0.0165 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.7990 0.1200 1.8490 0.5400 ;
        RECT 1.7990 0.5400 2.0940 0.5530 ;
        RECT 1.7990 0.5530 2.1830 0.5900 ;
        RECT 2.0440 0.5900 2.1830 0.6630 ;
        RECT 2.0440 0.6630 2.0940 0.7430 ;
        RECT 1.7990 0.7430 2.0940 0.7930 ;
        RECT 1.7990 0.7930 1.8490 1.5640 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Y
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 2.3950 1.7730 ;
    LAYER M1 ;
      RECT 1.5350 0.6400 1.9410 0.6900 ;
      RECT 1.5350 0.5110 1.5850 0.6400 ;
      RECT 1.5350 0.6900 1.5850 1.0210 ;
      RECT 1.4950 0.4610 1.5850 0.5110 ;
      RECT 1.4950 1.0210 1.5850 1.0710 ;
      RECT 1.4950 0.1200 1.5450 0.4610 ;
      RECT 1.4950 1.0710 1.5450 1.5640 ;
      RECT 0.9270 0.6720 1.1810 0.7060 ;
      RECT 0.8870 0.6560 1.1810 0.6720 ;
      RECT 0.8870 0.6220 0.9770 0.6560 ;
      RECT 0.2790 1.2630 0.9770 1.3130 ;
      RECT 0.8870 0.1210 0.9370 0.6220 ;
      RECT 0.8870 1.3130 0.9370 1.5590 ;
      RECT 0.9270 0.7060 0.9770 1.2630 ;
      RECT 0.5830 1.3130 0.6330 1.5590 ;
      RECT 0.2790 1.3130 0.3290 1.5590 ;
      RECT 1.2900 0.7290 1.4850 0.7790 ;
      RECT 1.2900 0.7790 1.3400 0.9400 ;
      RECT 1.2900 0.6010 1.3400 0.7290 ;
      RECT 1.1910 0.9400 1.3400 0.9900 ;
      RECT 1.1910 0.5530 1.3400 0.6010 ;
      RECT 1.1910 0.5510 1.3150 0.5530 ;
      RECT 1.1910 0.9900 1.2410 1.5570 ;
      RECT 1.1910 0.1170 1.2410 0.5510 ;
    LAYER PO ;
      RECT 1.2770 0.0720 1.3070 1.6090 ;
      RECT 1.4290 0.0620 1.4590 1.6090 ;
      RECT 1.1250 0.0720 1.1550 1.6090 ;
      RECT 0.9730 0.0710 1.0030 1.6090 ;
      RECT 0.6690 0.0710 0.6990 1.6090 ;
      RECT 0.3650 0.0710 0.3950 1.6090 ;
      RECT 0.5170 0.0710 0.5470 1.6090 ;
      RECT 0.2130 0.0710 0.2430 1.6090 ;
      RECT 0.8210 0.0710 0.8510 1.6090 ;
      RECT 0.0610 0.0710 0.0910 1.6090 ;
      RECT 1.7330 0.0620 1.7630 1.6090 ;
      RECT 1.8850 0.0620 1.9150 1.6090 ;
      RECT 2.1890 0.0620 2.2190 1.6090 ;
      RECT 2.0370 0.0620 2.0670 1.6090 ;
      RECT 1.5810 0.0620 1.6110 1.6090 ;
  END
END AND4X2_LVT

MACRO AND4X4_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.584 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 2.5840 1.7020 ;
        RECT 1.3430 0.8230 1.3930 1.6420 ;
        RECT 0.4310 1.3770 0.4810 1.6420 ;
        RECT 0.7350 1.3770 0.7850 1.6420 ;
        RECT 1.0390 1.1990 1.0890 1.6420 ;
        RECT 1.7990 1.0080 1.8490 1.6420 ;
        RECT 2.1030 1.0080 2.1530 1.6420 ;
    END
  END VDD

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 0.7350 0.7250 0.7850 ;
        RECT 0.5530 0.7050 0.6630 0.7350 ;
        RECT 0.5530 0.7850 0.6630 0.8150 ;
    END
    ANTENNAGATEAREA 0.0165 ;
  END A2

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7350 0.4210 0.7850 ;
        RECT 0.2490 0.7050 0.3590 0.7350 ;
        RECT 0.2490 0.7850 0.3590 0.8150 ;
    END
    ANTENNAGATEAREA 0.0165 ;
  END A4

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.6470 0.1150 1.6970 0.5140 ;
        RECT 1.6470 0.5140 2.4100 0.5530 ;
        RECT 1.9510 0.1150 2.0010 0.5140 ;
        RECT 2.2550 0.1150 2.3050 0.5140 ;
        RECT 1.6470 0.5530 2.4970 0.5640 ;
        RECT 2.3600 0.5640 2.4970 0.6630 ;
        RECT 2.3600 0.6630 2.4100 0.8260 ;
        RECT 1.6470 0.8260 2.4100 0.8760 ;
        RECT 1.6470 0.8760 1.6970 1.5650 ;
        RECT 1.9510 0.8760 2.0010 1.5650 ;
        RECT 2.2550 0.8760 2.3050 1.5650 ;
    END
    ANTENNADIFFAREA 0.3972 ;
  END Y

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 2.5840 0.0300 ;
        RECT 1.0390 0.0300 1.0890 0.3040 ;
        RECT 1.7990 0.0300 1.8490 0.4130 ;
        RECT 0.2790 0.0300 0.3290 0.4790 ;
        RECT 1.3430 0.0300 1.3930 0.4800 ;
        RECT 2.1030 0.0300 2.1530 0.4130 ;
    END
  END VSS

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 1.0090 0.5110 1.0390 ;
        RECT 0.4010 1.0390 0.5730 1.0890 ;
        RECT 0.4010 1.0890 0.5110 1.1190 ;
    END
    ANTENNAGATEAREA 0.0165 ;
  END A3

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 1.0090 0.8150 1.0390 ;
        RECT 0.7050 1.0390 0.8770 1.0890 ;
        RECT 0.7050 1.0890 0.8150 1.1190 ;
    END
    ANTENNAGATEAREA 0.0165 ;
  END A1
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 2.6990 1.7730 ;
    LAYER M1 ;
      RECT 0.8870 0.6560 1.1810 0.6720 ;
      RECT 0.9270 0.6720 1.1810 0.7060 ;
      RECT 0.8870 0.6220 0.9770 0.6560 ;
      RECT 0.8870 0.1210 0.9370 0.6220 ;
      RECT 0.2790 1.2630 0.9770 1.3130 ;
      RECT 0.8870 1.3130 0.9370 1.5590 ;
      RECT 0.9270 0.7060 0.9770 1.2630 ;
      RECT 0.5830 1.3130 0.6330 1.5590 ;
      RECT 0.2790 1.3130 0.3290 1.5590 ;
      RECT 1.5350 0.6420 2.2450 0.6920 ;
      RECT 1.5350 0.6920 1.5850 0.6980 ;
      RECT 1.5350 0.5050 1.5850 0.6420 ;
      RECT 1.4950 0.6980 1.5850 0.7480 ;
      RECT 1.4950 0.4550 1.5850 0.5050 ;
      RECT 1.4950 0.7480 1.5450 1.5640 ;
      RECT 1.4950 0.1140 1.5450 0.4550 ;
      RECT 1.2310 0.6010 1.4850 0.6490 ;
      RECT 1.1910 0.5990 1.4850 0.6010 ;
      RECT 1.2310 0.6490 1.2810 0.8720 ;
      RECT 1.1910 0.5510 1.2810 0.5990 ;
      RECT 1.1910 0.8720 1.2810 0.9220 ;
      RECT 1.1910 0.1170 1.2410 0.5510 ;
      RECT 1.1910 0.9220 1.2410 1.5570 ;
    LAYER PO ;
      RECT 0.0610 0.0710 0.0910 1.6090 ;
      RECT 0.8210 0.0710 0.8510 1.6090 ;
      RECT 0.2130 0.0710 0.2430 1.6090 ;
      RECT 0.5170 0.0710 0.5470 1.6090 ;
      RECT 0.3650 0.0710 0.3950 1.6090 ;
      RECT 0.6690 0.0710 0.6990 1.6090 ;
      RECT 0.9730 0.0710 1.0030 1.6090 ;
      RECT 1.1250 0.0720 1.1550 1.6090 ;
      RECT 1.4290 0.0640 1.4590 1.6170 ;
      RECT 1.2770 0.0720 1.3070 1.6090 ;
      RECT 1.5810 0.0640 1.6110 1.6080 ;
      RECT 1.8850 0.0720 1.9150 1.6100 ;
      RECT 2.0370 0.0720 2.0670 1.6100 ;
      RECT 2.1890 0.0720 2.2190 1.6100 ;
      RECT 2.4930 0.0720 2.5230 1.6100 ;
      RECT 2.3410 0.0720 2.3710 1.6100 ;
      RECT 1.7330 0.0720 1.7630 1.6100 ;
  END
END AND4X4_LVT

MACRO ANTENNA_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.456 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 0.4560 1.7020 ;
    END
  END VDD

  PIN INP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0970 0.7050 0.2560 0.8160 ;
        RECT 0.2000 0.8160 0.2560 1.1510 ;
        RECT 0.2000 0.2950 0.2560 0.7050 ;
    END
    ANTENNADIFFAREA 0.0805 ;
    ANTENNAGATEAREA 0.0805 ;
  END INP

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 0.4560 0.0300 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 0.5710 1.7730 ;
  END
END ANTENNA_LVT

MACRO AO21X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.52 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.5200 1.7020 ;
        RECT 0.5820 1.2050 0.6320 1.6420 ;
        RECT 0.2790 1.1130 0.3290 1.6420 ;
        RECT 1.0390 0.8280 1.0890 1.6420 ;
    END
  END VDD

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4920 0.8570 0.6630 0.9670 ;
    END
    ANTENNAGATEAREA 0.0243 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1610 1.1610 1.2710 1.2710 ;
        RECT 1.1910 1.2710 1.2410 1.5540 ;
        RECT 1.1910 0.8550 1.2410 1.1610 ;
        RECT 1.1910 0.8050 1.2810 0.8550 ;
        RECT 1.2310 0.4920 1.2810 0.8050 ;
        RECT 1.1910 0.4420 1.2810 0.4920 ;
        RECT 1.1910 0.1340 1.2410 0.4420 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.7050 0.4210 0.8150 ;
    END
    ANTENNAGATEAREA 0.0243 ;
  END A2

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.5200 0.0300 ;
        RECT 1.0400 0.0300 1.0900 0.4960 ;
        RECT 0.2790 0.0300 0.3290 0.2880 ;
        RECT 0.2790 0.2880 0.7850 0.3380 ;
        RECT 0.7350 0.3380 0.7850 0.5620 ;
        RECT 0.2790 0.3380 0.3290 0.5620 ;
    END
  END VSS

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 0.0970 0.8770 0.2070 ;
    END
    ANTENNAGATEAREA 0.0225 ;
  END A3
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.6350 1.7730 ;
    LAYER M1 ;
      RECT 0.5830 0.6200 1.1810 0.6700 ;
      RECT 0.5830 0.3880 0.6330 0.6200 ;
      RECT 0.8870 0.6700 0.9370 1.5680 ;
      RECT 0.8870 0.3880 0.9370 0.6200 ;
      RECT 0.7350 1.1200 0.7850 1.5630 ;
      RECT 0.4310 1.0700 0.7850 1.1200 ;
      RECT 0.4310 1.1200 0.4810 1.5680 ;
    LAYER PO ;
      RECT 1.2770 0.0630 1.3070 1.6040 ;
      RECT 0.2130 0.0640 0.2430 1.6130 ;
      RECT 1.1250 0.0640 1.1550 1.6040 ;
      RECT 0.8210 0.0590 0.8510 1.6130 ;
      RECT 0.9730 0.0640 1.0030 1.6130 ;
      RECT 0.6690 0.0640 0.6990 1.6130 ;
      RECT 0.0610 0.0640 0.0910 1.6130 ;
      RECT 1.4290 0.0630 1.4590 1.6040 ;
      RECT 0.3650 0.0590 0.3950 1.6130 ;
      RECT 0.5170 0.0640 0.5470 1.6130 ;
  END
END AO21X1_LVT

MACRO AO21X2_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.672 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3120 1.0090 1.4220 1.1190 ;
        RECT 1.3440 1.1190 1.3940 1.5440 ;
        RECT 1.3440 0.7500 1.3940 1.0090 ;
        RECT 1.3440 0.7000 1.4320 0.7500 ;
        RECT 1.3820 0.5180 1.4320 0.7000 ;
        RECT 1.0100 0.4680 1.4320 0.5180 ;
        RECT 1.3440 0.1600 1.3940 0.4680 ;
        RECT 1.0390 0.1600 1.0890 0.4680 ;
        RECT 1.0100 0.5180 1.0600 0.7440 ;
        RECT 1.0100 0.7440 1.0890 0.7940 ;
        RECT 1.0390 0.7940 1.0890 1.1020 ;
    END
    ANTENNADIFFAREA 0.2484 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4910 0.8570 0.6620 0.9670 ;
    END
    ANTENNAGATEAREA 0.0243 ;
  END A1

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.6720 0.0300 ;
        RECT 1.1910 0.0300 1.2410 0.3970 ;
        RECT 0.2790 0.0300 0.3290 0.2950 ;
        RECT 0.2790 0.2950 0.7850 0.3450 ;
        RECT 0.7350 0.3450 0.7850 0.5690 ;
        RECT 0.2790 0.3450 0.3290 0.5690 ;
    END
  END VSS

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2480 0.7050 0.4210 0.8150 ;
    END
    ANTENNAGATEAREA 0.0243 ;
  END A2

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.6720 1.7020 ;
        RECT 0.5830 1.2120 0.6330 1.6420 ;
        RECT 0.2790 1.1200 0.3290 1.6420 ;
        RECT 1.1910 1.2880 1.2410 1.6420 ;
    END
  END VDD

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7040 0.0970 0.8770 0.2070 ;
    END
    ANTENNAGATEAREA 0.0225 ;
  END A3
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.7870 1.7730 ;
    LAYER M1 ;
      RECT 1.1150 0.5680 1.3170 0.6500 ;
      RECT 1.1980 0.6500 1.2480 1.1520 ;
      RECT 0.8870 1.1520 1.2480 1.2020 ;
      RECT 0.5830 0.3950 0.6330 0.6510 ;
      RECT 0.8870 1.2020 0.9370 1.5750 ;
      RECT 0.8870 0.7010 0.9370 1.1520 ;
      RECT 0.5830 0.6510 0.9370 0.7010 ;
      RECT 0.8870 0.3950 0.9370 0.6510 ;
      RECT 0.7350 1.1270 0.7850 1.5700 ;
      RECT 0.4310 1.0770 0.7850 1.1270 ;
      RECT 0.4310 1.1270 0.4810 1.5750 ;
    LAYER PO ;
      RECT 1.4290 0.0560 1.4590 1.5970 ;
      RECT 0.5170 0.0710 0.5470 1.6200 ;
      RECT 1.5810 0.0560 1.6110 1.5970 ;
      RECT 0.0610 0.0640 0.0910 1.6130 ;
      RECT 0.6690 0.0710 0.6990 1.6200 ;
      RECT 0.3650 0.0660 0.3950 1.6200 ;
      RECT 0.8210 0.0660 0.8510 1.6200 ;
      RECT 1.2770 0.0520 1.3070 1.6040 ;
      RECT 0.9730 0.0640 1.0030 1.6130 ;
      RECT 1.1250 0.0640 1.1550 1.6040 ;
      RECT 0.2130 0.0640 0.2430 1.6130 ;
  END
END AO21X2_LVT

MACRO AO221X1_LVT
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.824 BY 1.672 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.0090 0.7730 1.1810 0.8230 ;
        RECT 1.0090 0.7050 1.1190 0.7730 ;
    END
    ANTENNAGATEAREA 0.021 ;
  END A5

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2490 0.8560 0.4040 0.9670 ;
        RECT 0.3540 0.8460 0.4040 0.8560 ;
    END
    ANTENNAGATEAREA 0.0249 ;
  END A1

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5530 1.0060 0.6630 1.1230 ;
        RECT 0.6130 0.9040 0.6630 1.0060 ;
        RECT 0.6130 0.8540 0.7250 0.9040 ;
    END
    ANTENNAGATEAREA 0.0249 ;
  END A4

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4650 1.1610 1.5750 1.2710 ;
        RECT 1.4950 1.2710 1.5450 1.5540 ;
        RECT 1.4950 0.8650 1.5450 1.1610 ;
        RECT 1.4950 0.8640 1.5850 0.8650 ;
        RECT 1.4950 0.8030 1.5950 0.8640 ;
        RECT 1.5450 0.5040 1.5950 0.8030 ;
        RECT 1.4950 0.4530 1.5950 0.5040 ;
        RECT 1.4950 0.1460 1.5450 0.4530 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0.0000 1.6420 1.8240 1.7020 ;
        RECT 0.4310 1.3740 0.4810 1.6420 ;
        RECT 1.3420 0.7350 1.3920 1.6420 ;
    END
  END VDD

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4010 0.5530 0.5730 0.6630 ;
    END
    ANTENNAGATEAREA 0.0249 ;
  END A2

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0.0000 -0.0300 1.8240 0.0300 ;
        RECT 1.0400 0.0300 1.0900 0.3660 ;
        RECT 0.5830 0.0300 0.6330 0.4710 ;
        RECT 1.3430 0.0300 1.3930 0.4840 ;
    END
  END VSS

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7050 0.0970 0.8630 0.2070 ;
    END
    ANTENNAGATEAREA 0.0249 ;
  END A3
  OBS
    LAYER NWELL ;
      RECT -0.1150 0.6790 1.9390 1.7730 ;
    LAYER M1 ;
      RECT 1.1910 0.6350 1.4850 0.6850 ;
      RECT 0.2790 0.2960 0.3290 0.7280 ;
      RECT 0.8870 0.5600 0.9370 0.7280 ;
      RECT 0.8870 0.3210 0.9370 0.5100 ;
      RECT 0.2790 0.7280 0.9370 0.7780 ;
      RECT 0.8870 0.7780 0.9370 0.9080 ;
      RECT 1.1910 0.5600 1.2410 0.6350 ;
      RECT 0.8870 0.5100 1.2410 0.5600 ;
      RECT 1.1910 0.2660 1.2410 0.5100 ;
      RECT 0.8870 0.9080 1.2410 0.9580 ;
      RECT 1.1910 0.9580 1.2410 1.5710 ;
      RECT 0.8870 1.3240 0.9370 1.5570 ;
      RECT 0.5830 1.3240 0.6330 1.5570 ;
      RECT 0.2790 1.2740 0.9370 1.3240 ;
      RECT 0.2790 1.3240 0.3290 1.5570 ;
      RECT 1.0390 1.0710 1.0890 1.5710 ;
      RECT 0.7350 1.0210 1.0890 1.0710 ;
      RECT 0.7350 1.0710 0.7850 1.2240 ;
    LAYER PO ;
      RECT 1.2770 0.0750 1.3070 1.6160 ;
      RECT 1.5810 0.0750 1.6110 1.6160 ;
      RECT 1.1250 0.0760 1.1550 1.6210 ;
      RECT 0.2130 0.0720 0.2430 1.6210 ;
      RECT 0.8210 0.0720 0.8510 1.6210 ;
      RECT 1.4290 0.0760 1.4590 1.6160 ;
      RECT 0.9730 0.0760 1.0030 1.6210 ;
      RECT 0.0610 0.0720 0.0910 1.6210 ;
      RECT 1.7330 0.0750 1.7630 1.6160 ;
      RECT 0.3650 0.0670 0.3950 1.6210 ;
      RECT 0.5170 0.0720 0.5470 1.6210 ;
      RECT 0.6690 0.0720 0.6990 1.6210 ;
  END
END AO221X1_LVT
  
END LIBRARY
